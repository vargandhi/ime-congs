module Queue_6_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 38515:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 38516:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 38517:4]
  output        io_enq_ready, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  input         io_enq_valid, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  input  [3:0]  io_enq_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  input  [31:0] io_enq_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  input  [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  input         io_deq_ready, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  output        io_deq_valid, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  output [3:0]  io_deq_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  output        io_deq_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  output [31:0] io_deq_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  output [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 38518:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  reg  ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  reg [31:0] ram_address [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [31:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38521:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38522:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 38523:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.RocketConfig.fir 38524:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.RocketConfig.fir 38525:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.RocketConfig.fir 38526:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.RocketConfig.fir 38527:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 38528:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 38531:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 38546:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 38552:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.RocketConfig.fir 38555:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  assign ram_param_MPORT_data = 3'h0;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  assign ram_source_MPORT_data = 1'h0;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.RocketConfig.fir 38561:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.RocketConfig.fir 38559:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38571:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38570:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38569:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38568:4]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38567:4]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38566:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38565:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38564:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38520:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38521:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38521:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.RocketConfig.fir 38534:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 38547:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38522:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38522:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.RocketConfig.fir 38549:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 38553:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 38523:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 38523:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.RocketConfig.fir 38556:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.RocketConfig.fir 38557:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_7_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 38579:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 38580:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 38581:4]
  output        io_enq_ready, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  input         io_enq_valid, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  input  [1:0]  io_enq_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  input  [3:0]  io_enq_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  input         io_enq_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  input  [2:0]  io_enq_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  input         io_enq_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  input         io_deq_ready, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  output        io_deq_valid, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  output [1:0]  io_deq_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  output [3:0]  io_deq_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  output        io_deq_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  output [2:0]  io_deq_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  output        io_deq_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 38582:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  reg  ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  reg [2:0] ram_sink [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire [2:0] ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire [2:0] ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38585:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38586:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 38587:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.RocketConfig.fir 38588:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.RocketConfig.fir 38589:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.RocketConfig.fir 38590:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.RocketConfig.fir 38591:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 38592:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 38595:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 38610:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 38616:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.RocketConfig.fir 38619:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_addr = value_1;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  assign ram_sink_MPORT_data = io_enq_bits_sink;
  assign ram_sink_MPORT_addr = value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.RocketConfig.fir 38625:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.RocketConfig.fir 38623:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38635:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38634:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38633:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38632:4]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38631:4]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38630:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38629:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 38628:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 38584:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38585:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38585:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.RocketConfig.fir 38598:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 38611:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38586:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 38586:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.RocketConfig.fir 38613:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 38617:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 38587:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 38587:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.RocketConfig.fir 38620:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.RocketConfig.fir 38621:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HellaPeekingArbiter_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 270408:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 270409:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 270410:4]
  output        io_in_1_ready, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input         io_in_1_valid, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [2:0]  io_in_1_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [2:0]  io_in_1_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [3:0]  io_in_1_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [3:0]  io_in_1_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [63:0] io_in_1_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input         io_in_1_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [7:0]  io_in_1_bits_union, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input         io_in_1_bits_last, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output        io_in_4_ready, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input         io_in_4_valid, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [2:0]  io_in_4_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [2:0]  io_in_4_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [3:0]  io_in_4_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [3:0]  io_in_4_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [31:0] io_in_4_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [63:0] io_in_4_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input         io_in_4_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input  [7:0]  io_in_4_bits_union, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input         io_in_4_bits_last, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  input         io_out_ready, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output        io_out_valid, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output [2:0]  io_out_bits_chanId, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output [2:0]  io_out_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output [2:0]  io_out_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output [3:0]  io_out_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output [3:0]  io_out_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output [31:0] io_out_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output [63:0] io_out_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output        io_out_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output [7:0]  io_out_bits_union, // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
  output        io_out_bits_last // @[chipyard.TestHarness.RocketConfig.fir 270411:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lockIdx; // @[Arbiters.scala 25:20 chipyard.TestHarness.RocketConfig.fir 270416:4]
  reg  locked; // @[Arbiters.scala 26:19 chipyard.TestHarness.RocketConfig.fir 270417:4]
  wire [2:0] choice = io_in_1_valid ? 3'h1 : 3'h4; // @[Mux.scala 47:69 chipyard.TestHarness.RocketConfig.fir 270420:4]
  wire [2:0] chosen = locked ? lockIdx : choice; // @[Arbiters.scala 36:19 chipyard.TestHarness.RocketConfig.fir 270422:4]
  wire  _io_in_1_ready_T = chosen == 3'h1; // @[Arbiters.scala 39:46 chipyard.TestHarness.RocketConfig.fir 270426:4]
  wire  _io_in_4_ready_T = chosen == 3'h4; // @[Arbiters.scala 39:46 chipyard.TestHarness.RocketConfig.fir 270435:4]
  wire [2:0] _GEN_14 = 3'h1 == chosen ? 3'h3 : 3'h4; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [2:0] _GEN_15 = 3'h1 == chosen ? io_in_1_bits_opcode : 3'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [2:0] _GEN_16 = 3'h1 == chosen ? io_in_1_bits_param : 3'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [3:0] _GEN_17 = 3'h1 == chosen ? io_in_1_bits_size : 4'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [3:0] _GEN_18 = 3'h1 == chosen ? io_in_1_bits_source : 4'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [63:0] _GEN_20 = 3'h1 == chosen ? io_in_1_bits_data : 64'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [7:0] _GEN_22 = 3'h1 == chosen ? io_in_1_bits_union : 8'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire  _GEN_23 = 3'h1 == chosen ? io_in_1_bits_last : 1'h1; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire  _GEN_25 = 3'h2 == chosen ? 1'h0 : 3'h1 == chosen & io_in_1_valid; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [2:0] _GEN_26 = 3'h2 == chosen ? 3'h2 : _GEN_14; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [2:0] _GEN_27 = 3'h2 == chosen ? 3'h0 : _GEN_15; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [2:0] _GEN_28 = 3'h2 == chosen ? 3'h0 : _GEN_16; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [3:0] _GEN_29 = 3'h2 == chosen ? 4'h0 : _GEN_17; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [3:0] _GEN_30 = 3'h2 == chosen ? 4'h0 : _GEN_18; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [63:0] _GEN_32 = 3'h2 == chosen ? 64'h0 : _GEN_20; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire  _GEN_33 = 3'h2 == chosen ? 1'h0 : 3'h1 == chosen & io_in_1_bits_corrupt; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [7:0] _GEN_34 = 3'h2 == chosen ? 8'h0 : _GEN_22; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire  _GEN_37 = 3'h3 == chosen ? 1'h0 : _GEN_25; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [2:0] _GEN_38 = 3'h3 == chosen ? 3'h1 : _GEN_26; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [2:0] _GEN_39 = 3'h3 == chosen ? 3'h0 : _GEN_27; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [2:0] _GEN_40 = 3'h3 == chosen ? 3'h0 : _GEN_28; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [3:0] _GEN_41 = 3'h3 == chosen ? 4'h0 : _GEN_29; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [3:0] _GEN_42 = 3'h3 == chosen ? 4'h0 : _GEN_30; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [63:0] _GEN_44 = 3'h3 == chosen ? 64'h0 : _GEN_32; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire  _GEN_45 = 3'h3 == chosen ? 1'h0 : _GEN_33; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire [7:0] _GEN_46 = 3'h3 == chosen ? 8'h0 : _GEN_34; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 270440:4]
  wire  _T_1 = ~locked; // @[Arbiters.scala 59:11 chipyard.TestHarness.RocketConfig.fir 270442:6]
  wire  _GEN_61 = _T_1 | locked; // @[Arbiters.scala 59:50 chipyard.TestHarness.RocketConfig.fir 270444:6 Arbiters.scala 61:14 chipyard.TestHarness.RocketConfig.fir 270446:8 Arbiters.scala 26:19 chipyard.TestHarness.RocketConfig.fir 270417:4]
  assign io_in_1_ready = io_out_ready & _io_in_1_ready_T; // @[Arbiters.scala 39:36 chipyard.TestHarness.RocketConfig.fir 270427:4]
  assign io_in_4_ready = io_out_ready & _io_in_4_ready_T; // @[Arbiters.scala 39:36 chipyard.TestHarness.RocketConfig.fir 270436:4]
  assign io_out_valid = 3'h4 == chosen ? io_in_4_valid : _GEN_37; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  assign io_out_bits_chanId = 3'h4 == chosen ? 3'h0 : _GEN_38; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  assign io_out_bits_opcode = 3'h4 == chosen ? io_in_4_bits_opcode : _GEN_39; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  assign io_out_bits_param = 3'h4 == chosen ? io_in_4_bits_param : _GEN_40; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  assign io_out_bits_size = 3'h4 == chosen ? io_in_4_bits_size : _GEN_41; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  assign io_out_bits_source = 3'h4 == chosen ? io_in_4_bits_source : _GEN_42; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  assign io_out_bits_address = 3'h4 == chosen ? io_in_4_bits_address : 32'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  assign io_out_bits_data = 3'h4 == chosen ? io_in_4_bits_data : _GEN_44; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  assign io_out_bits_corrupt = 3'h4 == chosen ? io_in_4_bits_corrupt : _GEN_45; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  assign io_out_bits_union = 3'h4 == chosen ? io_in_4_bits_union : _GEN_46; // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  assign io_out_bits_last = 3'h4 == chosen ? io_in_4_bits_last : 3'h3 == chosen | (3'h2 == chosen | _GEN_23); // @[Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4 Arbiters.scala 42:16 chipyard.TestHarness.RocketConfig.fir 270438:4]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiters.scala 25:20 chipyard.TestHarness.RocketConfig.fir 270416:4]
      lockIdx <= 3'h0; // @[Arbiters.scala 25:20 chipyard.TestHarness.RocketConfig.fir 270416:4]
    end else if (_T) begin // @[Arbiters.scala 58:24 chipyard.TestHarness.RocketConfig.fir 270441:4]
      if (_T_1) begin // @[Arbiters.scala 59:50 chipyard.TestHarness.RocketConfig.fir 270444:6]
        if (io_in_1_valid) begin // @[Mux.scala 47:69 chipyard.TestHarness.RocketConfig.fir 270420:4]
          lockIdx <= 3'h1;
        end else begin
          lockIdx <= 3'h4;
        end
      end
    end
    if (reset) begin // @[Arbiters.scala 26:19 chipyard.TestHarness.RocketConfig.fir 270417:4]
      locked <= 1'h0; // @[Arbiters.scala 26:19 chipyard.TestHarness.RocketConfig.fir 270417:4]
    end else if (_T) begin // @[Arbiters.scala 58:24 chipyard.TestHarness.RocketConfig.fir 270441:4]
      if (io_out_bits_last) begin // @[Arbiters.scala 64:35 chipyard.TestHarness.RocketConfig.fir 270448:6]
        locked <= 1'h0; // @[Arbiters.scala 65:14 chipyard.TestHarness.RocketConfig.fir 270449:8]
      end else begin
        locked <= _GEN_61;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockIdx = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  locked = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericSerializer_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 270453:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 270454:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 270455:4]
  output        io_in_ready, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input         io_in_valid, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input  [2:0]  io_in_bits_chanId, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input  [2:0]  io_in_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input  [2:0]  io_in_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input  [3:0]  io_in_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input  [3:0]  io_in_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input  [31:0] io_in_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input  [63:0] io_in_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input         io_in_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input  [7:0]  io_in_bits_union, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input         io_in_bits_last, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  input         io_out_ready, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  output        io_out_valid, // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
  output [3:0]  io_out_bits // @[chipyard.TestHarness.RocketConfig.fir 270456:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [122:0] data; // @[Serdes.scala 175:17 chipyard.TestHarness.RocketConfig.fir 270458:4]
  reg  sending; // @[Serdes.scala 177:24 chipyard.TestHarness.RocketConfig.fir 270459:4]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 270460:4]
  reg [4:0] sendCount; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 270461:4]
  wire  wrap_wrap = sendCount == 5'h1e; // @[Counter.scala 72:24 chipyard.TestHarness.RocketConfig.fir 270465:6]
  wire [4:0] _wrap_value_T_1 = sendCount + 5'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 270467:6]
  wire  sendDone = _T & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 270464:4 Counter.scala 118:24 chipyard.TestHarness.RocketConfig.fir 270472:6 chipyard.TestHarness.RocketConfig.fir 270463:4]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 270479:4]
  wire [122:0] _data_T = {io_in_bits_chanId,io_in_bits_opcode,io_in_bits_param,io_in_bits_size,io_in_bits_source,
    io_in_bits_address,io_in_bits_data,io_in_bits_corrupt,io_in_bits_union,io_in_bits_last}; // @[Serdes.scala 185:24 chipyard.TestHarness.RocketConfig.fir 270489:6]
  wire  _GEN_4 = _T_1 | sending; // @[Serdes.scala 184:23 chipyard.TestHarness.RocketConfig.fir 270480:4 Serdes.scala 186:13 chipyard.TestHarness.RocketConfig.fir 270491:6 Serdes.scala 177:24 chipyard.TestHarness.RocketConfig.fir 270459:4]
  wire [122:0] _data_T_1 = {{4'd0}, data[122:4]}; // @[Serdes.scala 189:39 chipyard.TestHarness.RocketConfig.fir 270495:6]
  assign io_in_ready = ~sending; // @[Serdes.scala 180:18 chipyard.TestHarness.RocketConfig.fir 270474:4]
  assign io_out_valid = sending; // @[Serdes.scala 181:16 chipyard.TestHarness.RocketConfig.fir 270476:4]
  assign io_out_bits = data[3:0]; // @[Serdes.scala 182:22 chipyard.TestHarness.RocketConfig.fir 270477:4]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 189:24 chipyard.TestHarness.RocketConfig.fir 270494:4]
      data <= _data_T_1; // @[Serdes.scala 189:31 chipyard.TestHarness.RocketConfig.fir 270496:6]
    end else if (_T_1) begin // @[Serdes.scala 184:23 chipyard.TestHarness.RocketConfig.fir 270480:4]
      data <= _data_T; // @[Serdes.scala 185:10 chipyard.TestHarness.RocketConfig.fir 270490:6]
    end
    if (reset) begin // @[Serdes.scala 177:24 chipyard.TestHarness.RocketConfig.fir 270459:4]
      sending <= 1'h0; // @[Serdes.scala 177:24 chipyard.TestHarness.RocketConfig.fir 270459:4]
    end else if (sendDone) begin // @[Serdes.scala 191:19 chipyard.TestHarness.RocketConfig.fir 270498:4]
      sending <= 1'h0; // @[Serdes.scala 191:29 chipyard.TestHarness.RocketConfig.fir 270499:6]
    end else begin
      sending <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 270461:4]
      sendCount <= 5'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 270461:4]
    end else if (_T) begin // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 270464:4]
      if (wrap_wrap) begin // @[Counter.scala 86:20 chipyard.TestHarness.RocketConfig.fir 270469:6]
        sendCount <= 5'h0; // @[Counter.scala 86:28 chipyard.TestHarness.RocketConfig.fir 270470:8]
      end else begin
        sendCount <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 270468:6]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  data = _RAND_0[122:0];
  _RAND_1 = {1{`RANDOM}};
  sending = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sendCount = _RAND_2[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericDeserializer_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 270502:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 270503:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 270504:4]
  output        io_in_ready, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  input         io_in_valid, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  input  [3:0]  io_in_bits, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  input         io_out_ready, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  output        io_out_valid, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  output [2:0]  io_out_bits_chanId, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  output [2:0]  io_out_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  output [2:0]  io_out_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  output [3:0]  io_out_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  output [3:0]  io_out_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  output [31:0] io_out_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  output [63:0] io_out_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  output        io_out_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
  output [7:0]  io_out_bits_union // @[chipyard.TestHarness.RocketConfig.fir 270505:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] data_0; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_1; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_2; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_3; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_4; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_5; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_6; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_7; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_8; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_9; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_10; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_11; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_12; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_13; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_14; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_15; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_16; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_17; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_18; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_19; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_20; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_21; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_22; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_23; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_24; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_25; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_26; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_27; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_28; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_29; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg [3:0] data_30; // @[Serdes.scala 202:17 chipyard.TestHarness.RocketConfig.fir 270507:4]
  reg  receiving; // @[Serdes.scala 204:26 chipyard.TestHarness.RocketConfig.fir 270508:4]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 270509:4]
  reg [4:0] recvCount; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 270510:4]
  wire  wrap_wrap = recvCount == 5'h1e; // @[Counter.scala 72:24 chipyard.TestHarness.RocketConfig.fir 270514:6]
  wire [4:0] _wrap_value_T_1 = recvCount + 5'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 270516:6]
  wire  recvDone = _T & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 270513:4 Counter.scala 118:24 chipyard.TestHarness.RocketConfig.fir 270521:6 chipyard.TestHarness.RocketConfig.fir 270512:4]
  wire [27:0] io_out_bits_lo_lo = {data_6,data_5,data_4,data_3,data_2,data_1,data_0}; // @[Serdes.scala 209:23 chipyard.TestHarness.RocketConfig.fir 270531:4]
  wire [59:0] io_out_bits_lo = {data_14,data_13,data_12,data_11,data_10,data_9,data_8,data_7,io_out_bits_lo_lo}; // @[Serdes.scala 209:23 chipyard.TestHarness.RocketConfig.fir 270539:4]
  wire [31:0] io_out_bits_hi_lo = {data_22,data_21,data_20,data_19,data_18,data_17,data_16,data_15}; // @[Serdes.scala 209:23 chipyard.TestHarness.RocketConfig.fir 270546:4]
  wire [123:0] _io_out_bits_T = {data_30,data_29,data_28,data_27,data_26,data_25,data_24,data_23,io_out_bits_hi_lo,
    io_out_bits_lo}; // @[Serdes.scala 209:23 chipyard.TestHarness.RocketConfig.fir 270555:4]
  wire  _GEN_65 = recvDone ? 1'h0 : receiving; // @[Serdes.scala 215:19 chipyard.TestHarness.RocketConfig.fir 270593:4 Serdes.scala 215:31 chipyard.TestHarness.RocketConfig.fir 270594:6 Serdes.scala 204:26 chipyard.TestHarness.RocketConfig.fir 270508:4]
  wire  _T_2 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 270596:4]
  wire  _GEN_66 = _T_2 | _GEN_65; // @[Serdes.scala 217:24 chipyard.TestHarness.RocketConfig.fir 270597:4 Serdes.scala 217:36 chipyard.TestHarness.RocketConfig.fir 270598:6]
  assign io_in_ready = receiving; // @[Serdes.scala 207:15 chipyard.TestHarness.RocketConfig.fir 270523:4]
  assign io_out_valid = ~receiving; // @[Serdes.scala 208:19 chipyard.TestHarness.RocketConfig.fir 270524:4]
  assign io_out_bits_chanId = _io_out_bits_T[122:120]; // @[Serdes.scala 209:38 chipyard.TestHarness.RocketConfig.fir 270577:4]
  assign io_out_bits_opcode = _io_out_bits_T[119:117]; // @[Serdes.scala 209:38 chipyard.TestHarness.RocketConfig.fir 270575:4]
  assign io_out_bits_param = _io_out_bits_T[116:114]; // @[Serdes.scala 209:38 chipyard.TestHarness.RocketConfig.fir 270573:4]
  assign io_out_bits_size = _io_out_bits_T[113:110]; // @[Serdes.scala 209:38 chipyard.TestHarness.RocketConfig.fir 270571:4]
  assign io_out_bits_source = _io_out_bits_T[109:106]; // @[Serdes.scala 209:38 chipyard.TestHarness.RocketConfig.fir 270569:4]
  assign io_out_bits_address = _io_out_bits_T[105:74]; // @[Serdes.scala 209:38 chipyard.TestHarness.RocketConfig.fir 270567:4]
  assign io_out_bits_data = _io_out_bits_T[73:10]; // @[Serdes.scala 209:38 chipyard.TestHarness.RocketConfig.fir 270565:4]
  assign io_out_bits_corrupt = _io_out_bits_T[9]; // @[Serdes.scala 209:38 chipyard.TestHarness.RocketConfig.fir 270563:4]
  assign io_out_bits_union = _io_out_bits_T[8:1]; // @[Serdes.scala 209:38 chipyard.TestHarness.RocketConfig.fir 270561:4]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h0 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_0 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h1 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_1 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h2 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_2 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h3 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_3 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h4 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_4 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h5 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_5 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h6 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_6 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h7 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_7 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h8 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_8 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h9 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_9 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'ha == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_10 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'hb == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_11 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'hc == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_12 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'hd == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_13 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'he == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_14 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'hf == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_15 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h10 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_16 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h11 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_17 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h12 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_18 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h13 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_19 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h14 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_20 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h15 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_21 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h16 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_22 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h17 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_23 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h18 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_24 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h19 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_25 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h1a == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_26 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h1b == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_27 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h1c == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_28 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h1d == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_29 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.RocketConfig.fir 270590:4]
      if (5'h1e == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
        data_30 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.RocketConfig.fir 270591:6]
      end
    end
    receiving <= reset | _GEN_66; // @[Serdes.scala 204:26 chipyard.TestHarness.RocketConfig.fir 270508:4 Serdes.scala 204:26 chipyard.TestHarness.RocketConfig.fir 270508:4]
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 270510:4]
      recvCount <= 5'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 270510:4]
    end else if (_T) begin // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 270513:4]
      if (wrap_wrap) begin // @[Counter.scala 86:20 chipyard.TestHarness.RocketConfig.fir 270518:6]
        recvCount <= 5'h0; // @[Counter.scala 86:28 chipyard.TestHarness.RocketConfig.fir 270519:8]
      end else begin
        recvCount <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 270517:6]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  data_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  data_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  data_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  data_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  data_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  data_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  data_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  data_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  data_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  data_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  data_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  data_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  data_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  data_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  data_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  data_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  data_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  data_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  data_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  data_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  data_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  data_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  data_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  data_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  data_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  data_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  data_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  data_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  data_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  data_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  receiving = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  recvCount = _RAND_32[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SerialAdapter_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 281578:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 281579:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 281580:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 281581:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 281581:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 281581:4]
  output [3:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 281581:4]
  output [31:0] auto_out_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 281581:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 281581:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 281581:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 281581:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 281581:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 281581:4]
  output        io_serial_in_ready, // @[chipyard.TestHarness.RocketConfig.fir 281582:4]
  input         io_serial_in_valid, // @[chipyard.TestHarness.RocketConfig.fir 281582:4]
  input  [31:0] io_serial_in_bits, // @[chipyard.TestHarness.RocketConfig.fir 281582:4]
  input         io_serial_out_ready, // @[chipyard.TestHarness.RocketConfig.fir 281582:4]
  output        io_serial_out_valid, // @[chipyard.TestHarness.RocketConfig.fir 281582:4]
  output [31:0] io_serial_out_bits // @[chipyard.TestHarness.RocketConfig.fir 281582:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cmd; // @[SerialAdapter.scala 86:16 chipyard.TestHarness.RocketConfig.fir 281591:4]
  reg [63:0] addr; // @[SerialAdapter.scala 87:17 chipyard.TestHarness.RocketConfig.fir 281592:4]
  reg [63:0] len; // @[SerialAdapter.scala 88:16 chipyard.TestHarness.RocketConfig.fir 281593:4]
  reg [31:0] body_0; // @[SerialAdapter.scala 89:17 chipyard.TestHarness.RocketConfig.fir 281594:4]
  reg [31:0] body_1; // @[SerialAdapter.scala 89:17 chipyard.TestHarness.RocketConfig.fir 281594:4]
  reg [1:0] bodyValid; // @[SerialAdapter.scala 90:22 chipyard.TestHarness.RocketConfig.fir 281595:4]
  reg  idx; // @[SerialAdapter.scala 91:16 chipyard.TestHarness.RocketConfig.fir 281596:4]
  reg [3:0] state; // @[SerialAdapter.scala 97:22 chipyard.TestHarness.RocketConfig.fir 281597:4]
  wire  _io_serial_in_ready_T = state == 4'h0; // @[package.scala 15:47 chipyard.TestHarness.RocketConfig.fir 281598:4]
  wire  _io_serial_in_ready_T_1 = state == 4'h1; // @[package.scala 15:47 chipyard.TestHarness.RocketConfig.fir 281599:4]
  wire  _io_serial_in_ready_T_2 = state == 4'h2; // @[package.scala 15:47 chipyard.TestHarness.RocketConfig.fir 281600:4]
  wire  _io_serial_in_ready_T_3 = state == 4'h6; // @[package.scala 15:47 chipyard.TestHarness.RocketConfig.fir 281601:4]
  wire  _io_serial_in_ready_T_4 = _io_serial_in_ready_T | _io_serial_in_ready_T_1; // @[package.scala 72:59 chipyard.TestHarness.RocketConfig.fir 281602:4]
  wire  _io_serial_in_ready_T_5 = _io_serial_in_ready_T_4 | _io_serial_in_ready_T_2; // @[package.scala 72:59 chipyard.TestHarness.RocketConfig.fir 281603:4]
  wire  _io_serial_out_valid_T = state == 4'h5; // @[SerialAdapter.scala 100:32 chipyard.TestHarness.RocketConfig.fir 281606:4]
  wire [28:0] beatAddr = addr[31:3]; // @[SerialAdapter.scala 103:22 chipyard.TestHarness.RocketConfig.fir 281609:4]
  wire [28:0] nextAddr_hi = beatAddr + 29'h1; // @[SerialAdapter.scala 104:31 chipyard.TestHarness.RocketConfig.fir 281611:4]
  wire [31:0] nextAddr = {nextAddr_hi,3'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 281612:4]
  wire [3:0] wmask_lo = bodyValid[0] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12 chipyard.TestHarness.RocketConfig.fir 281616:4]
  wire [3:0] wmask_hi = bodyValid[1] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12 chipyard.TestHarness.RocketConfig.fir 281618:4]
  wire [7:0] wmask = {wmask_hi,wmask_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 281619:4]
  wire [63:0] _GEN_55 = {{32'd0}, nextAddr}; // @[SerialAdapter.scala 107:28 chipyard.TestHarness.RocketConfig.fir 281620:4]
  wire [63:0] addr_size = _GEN_55 - addr; // @[SerialAdapter.scala 107:28 chipyard.TestHarness.RocketConfig.fir 281621:4]
  wire [63:0] len_size_hi = len + 64'h1; // @[SerialAdapter.scala 108:26 chipyard.TestHarness.RocketConfig.fir 281623:4]
  wire [65:0] len_size = {len_size_hi,2'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 281624:4]
  wire [65:0] _GEN_56 = {{2'd0}, addr_size}; // @[SerialAdapter.scala 109:31 chipyard.TestHarness.RocketConfig.fir 281625:4]
  wire  _raw_size_T = len_size < _GEN_56; // @[SerialAdapter.scala 109:31 chipyard.TestHarness.RocketConfig.fir 281625:4]
  wire [65:0] raw_size = _raw_size_T ? len_size : {{2'd0}, addr_size}; // @[SerialAdapter.scala 109:21 chipyard.TestHarness.RocketConfig.fir 281626:4]
  wire  _rsize_T = 66'h1 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.RocketConfig.fir 281627:4]
  wire [1:0] _rsize_T_1 = _rsize_T ? 2'h0 : 2'h3; // @[Mux.scala 80:57 chipyard.TestHarness.RocketConfig.fir 281628:4]
  wire  _rsize_T_2 = 66'h2 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.RocketConfig.fir 281629:4]
  wire [1:0] _rsize_T_3 = _rsize_T_2 ? 2'h1 : _rsize_T_1; // @[Mux.scala 80:57 chipyard.TestHarness.RocketConfig.fir 281630:4]
  wire  _rsize_T_4 = 66'h4 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.RocketConfig.fir 281631:4]
  wire [1:0] rsize = _rsize_T_4 ? 2'h2 : _rsize_T_3; // @[Mux.scala 80:57 chipyard.TestHarness.RocketConfig.fir 281632:4]
  wire [1:0] _pow2size_T_66 = raw_size[0] + raw_size[1]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281699:4]
  wire [1:0] _pow2size_T_68 = raw_size[2] + raw_size[3]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281701:4]
  wire [2:0] _pow2size_T_70 = _pow2size_T_66 + _pow2size_T_68; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281703:4]
  wire [1:0] _pow2size_T_72 = raw_size[4] + raw_size[5]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281705:4]
  wire [1:0] _pow2size_T_74 = raw_size[6] + raw_size[7]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281707:4]
  wire [2:0] _pow2size_T_76 = _pow2size_T_72 + _pow2size_T_74; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281709:4]
  wire [3:0] _pow2size_T_78 = _pow2size_T_70 + _pow2size_T_76; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281711:4]
  wire [1:0] _pow2size_T_80 = raw_size[8] + raw_size[9]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281713:4]
  wire [1:0] _pow2size_T_82 = raw_size[10] + raw_size[11]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281715:4]
  wire [2:0] _pow2size_T_84 = _pow2size_T_80 + _pow2size_T_82; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281717:4]
  wire [1:0] _pow2size_T_86 = raw_size[12] + raw_size[13]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281719:4]
  wire [1:0] _pow2size_T_88 = raw_size[14] + raw_size[15]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281721:4]
  wire [2:0] _pow2size_T_90 = _pow2size_T_86 + _pow2size_T_88; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281723:4]
  wire [3:0] _pow2size_T_92 = _pow2size_T_84 + _pow2size_T_90; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281725:4]
  wire [4:0] _pow2size_T_94 = _pow2size_T_78 + _pow2size_T_92; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281727:4]
  wire [1:0] _pow2size_T_96 = raw_size[16] + raw_size[17]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281729:4]
  wire [1:0] _pow2size_T_98 = raw_size[18] + raw_size[19]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281731:4]
  wire [2:0] _pow2size_T_100 = _pow2size_T_96 + _pow2size_T_98; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281733:4]
  wire [1:0] _pow2size_T_102 = raw_size[20] + raw_size[21]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281735:4]
  wire [1:0] _pow2size_T_104 = raw_size[22] + raw_size[23]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281737:4]
  wire [2:0] _pow2size_T_106 = _pow2size_T_102 + _pow2size_T_104; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281739:4]
  wire [3:0] _pow2size_T_108 = _pow2size_T_100 + _pow2size_T_106; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281741:4]
  wire [1:0] _pow2size_T_110 = raw_size[24] + raw_size[25]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281743:4]
  wire [1:0] _pow2size_T_112 = raw_size[26] + raw_size[27]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281745:4]
  wire [2:0] _pow2size_T_114 = _pow2size_T_110 + _pow2size_T_112; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281747:4]
  wire [1:0] _pow2size_T_116 = raw_size[28] + raw_size[29]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281749:4]
  wire [1:0] _pow2size_T_118 = raw_size[31] + raw_size[32]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281751:4]
  wire [1:0] _GEN_57 = {{1'd0}, raw_size[30]}; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281753:4]
  wire [2:0] _pow2size_T_120 = _GEN_57 + _pow2size_T_118; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281753:4]
  wire [2:0] _pow2size_T_122 = _pow2size_T_116 + _pow2size_T_120[1:0]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281755:4]
  wire [3:0] _pow2size_T_124 = _pow2size_T_114 + _pow2size_T_122; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281757:4]
  wire [4:0] _pow2size_T_126 = _pow2size_T_108 + _pow2size_T_124; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281759:4]
  wire [5:0] _pow2size_T_128 = _pow2size_T_94 + _pow2size_T_126; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281761:4]
  wire [1:0] _pow2size_T_130 = raw_size[33] + raw_size[34]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281763:4]
  wire [1:0] _pow2size_T_132 = raw_size[35] + raw_size[36]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281765:4]
  wire [2:0] _pow2size_T_134 = _pow2size_T_130 + _pow2size_T_132; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281767:4]
  wire [1:0] _pow2size_T_136 = raw_size[37] + raw_size[38]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281769:4]
  wire [1:0] _pow2size_T_138 = raw_size[39] + raw_size[40]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281771:4]
  wire [2:0] _pow2size_T_140 = _pow2size_T_136 + _pow2size_T_138; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281773:4]
  wire [3:0] _pow2size_T_142 = _pow2size_T_134 + _pow2size_T_140; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281775:4]
  wire [1:0] _pow2size_T_144 = raw_size[41] + raw_size[42]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281777:4]
  wire [1:0] _pow2size_T_146 = raw_size[43] + raw_size[44]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281779:4]
  wire [2:0] _pow2size_T_148 = _pow2size_T_144 + _pow2size_T_146; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281781:4]
  wire [1:0] _pow2size_T_150 = raw_size[45] + raw_size[46]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281783:4]
  wire [1:0] _pow2size_T_152 = raw_size[47] + raw_size[48]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281785:4]
  wire [2:0] _pow2size_T_154 = _pow2size_T_150 + _pow2size_T_152; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281787:4]
  wire [3:0] _pow2size_T_156 = _pow2size_T_148 + _pow2size_T_154; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281789:4]
  wire [4:0] _pow2size_T_158 = _pow2size_T_142 + _pow2size_T_156; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281791:4]
  wire [1:0] _pow2size_T_160 = raw_size[49] + raw_size[50]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281793:4]
  wire [1:0] _pow2size_T_162 = raw_size[51] + raw_size[52]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281795:4]
  wire [2:0] _pow2size_T_164 = _pow2size_T_160 + _pow2size_T_162; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281797:4]
  wire [1:0] _pow2size_T_166 = raw_size[53] + raw_size[54]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281799:4]
  wire [1:0] _pow2size_T_168 = raw_size[55] + raw_size[56]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281801:4]
  wire [2:0] _pow2size_T_170 = _pow2size_T_166 + _pow2size_T_168; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281803:4]
  wire [3:0] _pow2size_T_172 = _pow2size_T_164 + _pow2size_T_170; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281805:4]
  wire [1:0] _pow2size_T_174 = raw_size[57] + raw_size[58]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281807:4]
  wire [1:0] _pow2size_T_176 = raw_size[59] + raw_size[60]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281809:4]
  wire [2:0] _pow2size_T_178 = _pow2size_T_174 + _pow2size_T_176; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281811:4]
  wire [1:0] _pow2size_T_180 = raw_size[61] + raw_size[62]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281813:4]
  wire [1:0] _pow2size_T_182 = raw_size[64] + raw_size[65]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281815:4]
  wire [1:0] _GEN_58 = {{1'd0}, raw_size[63]}; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281817:4]
  wire [2:0] _pow2size_T_184 = _GEN_58 + _pow2size_T_182; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281817:4]
  wire [2:0] _pow2size_T_186 = _pow2size_T_180 + _pow2size_T_184[1:0]; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281819:4]
  wire [3:0] _pow2size_T_188 = _pow2size_T_178 + _pow2size_T_186; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281821:4]
  wire [4:0] _pow2size_T_190 = _pow2size_T_172 + _pow2size_T_188; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281823:4]
  wire [5:0] _pow2size_T_192 = _pow2size_T_158 + _pow2size_T_190; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281825:4]
  wire [6:0] _pow2size_T_194 = _pow2size_T_128 + _pow2size_T_192; // @[Bitwise.scala 47:55 chipyard.TestHarness.RocketConfig.fir 281827:4]
  wire  pow2size = _pow2size_T_194 == 7'h1; // @[SerialAdapter.scala 113:37 chipyard.TestHarness.RocketConfig.fir 281829:4]
  wire [2:0] byteAddr = pow2size ? addr[2:0] : 3'h0; // @[SerialAdapter.scala 114:21 chipyard.TestHarness.RocketConfig.fir 281831:4]
  wire [31:0] put_acquire_address = {beatAddr, 3'h0}; // @[SerialAdapter.scala 117:19 chipyard.TestHarness.RocketConfig.fir 281832:4]
  wire [63:0] put_acquire_data = {body_1,body_0}; // @[SerialAdapter.scala 118:10 chipyard.TestHarness.RocketConfig.fir 281833:4]
  wire [31:0] get_acquire_address = {beatAddr,byteAddr}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 281898:4]
  wire [2:0] _get_acquire_a_mask_sizeOH_T = {{1'd0}, rsize}; // @[Misc.scala 201:34 chipyard.TestHarness.RocketConfig.fir 281964:4]
  wire [1:0] get_acquire_a_mask_sizeOH_shiftAmount = _get_acquire_a_mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.RocketConfig.fir 281965:4]
  wire [3:0] _get_acquire_a_mask_sizeOH_T_1 = 4'h1 << get_acquire_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.RocketConfig.fir 281966:4]
  wire [2:0] get_acquire_a_mask_sizeOH = _get_acquire_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.RocketConfig.fir 281968:4]
  wire  _get_acquire_a_mask_T = rsize >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.RocketConfig.fir 281969:4]
  wire  get_acquire_a_mask_size = get_acquire_a_mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 281970:4]
  wire  get_acquire_a_mask_bit = get_acquire_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 281971:4]
  wire  get_acquire_a_mask_nbit = ~get_acquire_a_mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 281972:4]
  wire  _get_acquire_a_mask_acc_T = get_acquire_a_mask_size & get_acquire_a_mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 281974:4]
  wire  get_acquire_a_mask_acc = _get_acquire_a_mask_T | _get_acquire_a_mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 281975:4]
  wire  _get_acquire_a_mask_acc_T_1 = get_acquire_a_mask_size & get_acquire_a_mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 281977:4]
  wire  get_acquire_a_mask_acc_1 = _get_acquire_a_mask_T | _get_acquire_a_mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 281978:4]
  wire  get_acquire_a_mask_size_1 = get_acquire_a_mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 281979:4]
  wire  get_acquire_a_mask_bit_1 = get_acquire_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 281980:4]
  wire  get_acquire_a_mask_nbit_1 = ~get_acquire_a_mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 281981:4]
  wire  get_acquire_a_mask_eq_2 = get_acquire_a_mask_nbit & get_acquire_a_mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 281982:4]
  wire  _get_acquire_a_mask_acc_T_2 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 281983:4]
  wire  get_acquire_a_mask_acc_2 = get_acquire_a_mask_acc | _get_acquire_a_mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 281984:4]
  wire  get_acquire_a_mask_eq_3 = get_acquire_a_mask_nbit & get_acquire_a_mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 281985:4]
  wire  _get_acquire_a_mask_acc_T_3 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 281986:4]
  wire  get_acquire_a_mask_acc_3 = get_acquire_a_mask_acc | _get_acquire_a_mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 281987:4]
  wire  get_acquire_a_mask_eq_4 = get_acquire_a_mask_bit & get_acquire_a_mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 281988:4]
  wire  _get_acquire_a_mask_acc_T_4 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 281989:4]
  wire  get_acquire_a_mask_acc_4 = get_acquire_a_mask_acc_1 | _get_acquire_a_mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 281990:4]
  wire  get_acquire_a_mask_eq_5 = get_acquire_a_mask_bit & get_acquire_a_mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 281991:4]
  wire  _get_acquire_a_mask_acc_T_5 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 281992:4]
  wire  get_acquire_a_mask_acc_5 = get_acquire_a_mask_acc_1 | _get_acquire_a_mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 281993:4]
  wire  get_acquire_a_mask_size_2 = get_acquire_a_mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 281994:4]
  wire  get_acquire_a_mask_bit_2 = get_acquire_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 281995:4]
  wire  get_acquire_a_mask_nbit_2 = ~get_acquire_a_mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 281996:4]
  wire  get_acquire_a_mask_eq_6 = get_acquire_a_mask_eq_2 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 281997:4]
  wire  _get_acquire_a_mask_acc_T_6 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 281998:4]
  wire  get_acquire_a_mask_lo_lo_lo = get_acquire_a_mask_acc_2 | _get_acquire_a_mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 281999:4]
  wire  get_acquire_a_mask_eq_7 = get_acquire_a_mask_eq_2 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282000:4]
  wire  _get_acquire_a_mask_acc_T_7 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282001:4]
  wire  get_acquire_a_mask_lo_lo_hi = get_acquire_a_mask_acc_2 | _get_acquire_a_mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282002:4]
  wire  get_acquire_a_mask_eq_8 = get_acquire_a_mask_eq_3 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282003:4]
  wire  _get_acquire_a_mask_acc_T_8 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282004:4]
  wire  get_acquire_a_mask_lo_hi_lo = get_acquire_a_mask_acc_3 | _get_acquire_a_mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282005:4]
  wire  get_acquire_a_mask_eq_9 = get_acquire_a_mask_eq_3 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282006:4]
  wire  _get_acquire_a_mask_acc_T_9 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282007:4]
  wire  get_acquire_a_mask_lo_hi_hi = get_acquire_a_mask_acc_3 | _get_acquire_a_mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282008:4]
  wire  get_acquire_a_mask_eq_10 = get_acquire_a_mask_eq_4 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282009:4]
  wire  _get_acquire_a_mask_acc_T_10 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282010:4]
  wire  get_acquire_a_mask_hi_lo_lo = get_acquire_a_mask_acc_4 | _get_acquire_a_mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282011:4]
  wire  get_acquire_a_mask_eq_11 = get_acquire_a_mask_eq_4 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282012:4]
  wire  _get_acquire_a_mask_acc_T_11 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282013:4]
  wire  get_acquire_a_mask_hi_lo_hi = get_acquire_a_mask_acc_4 | _get_acquire_a_mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282014:4]
  wire  get_acquire_a_mask_eq_12 = get_acquire_a_mask_eq_5 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282015:4]
  wire  _get_acquire_a_mask_acc_T_12 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282016:4]
  wire  get_acquire_a_mask_hi_hi_lo = get_acquire_a_mask_acc_5 | _get_acquire_a_mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282017:4]
  wire  get_acquire_a_mask_eq_13 = get_acquire_a_mask_eq_5 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282018:4]
  wire  _get_acquire_a_mask_acc_T_13 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282019:4]
  wire  get_acquire_a_mask_hi_hi_hi = get_acquire_a_mask_acc_5 | _get_acquire_a_mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282020:4]
  wire [7:0] get_acquire_mask = {get_acquire_a_mask_hi_hi_hi,get_acquire_a_mask_hi_hi_lo,get_acquire_a_mask_hi_lo_hi,
    get_acquire_a_mask_hi_lo_lo,get_acquire_a_mask_lo_hi_hi,get_acquire_a_mask_lo_hi_lo,get_acquire_a_mask_lo_lo_hi,
    get_acquire_a_mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 282027:4]
  wire  _bundleOut_0_a_valid_T = state == 4'h7; // @[package.scala 15:47 chipyard.TestHarness.RocketConfig.fir 282031:4]
  wire  _bundleOut_0_a_valid_T_1 = state == 4'h3; // @[package.scala 15:47 chipyard.TestHarness.RocketConfig.fir 282032:4]
  wire [3:0] get_acquire_size = {{2'd0}, rsize}; // @[Edges.scala 447:17 chipyard.TestHarness.RocketConfig.fir 281957:4 Edges.scala 450:15 chipyard.TestHarness.RocketConfig.fir 281961:4]
  wire  _bundleOut_0_d_ready_T = state == 4'h8; // @[package.scala 15:47 chipyard.TestHarness.RocketConfig.fir 282051:4]
  wire  _bundleOut_0_d_ready_T_1 = state == 4'h4; // @[package.scala 15:47 chipyard.TestHarness.RocketConfig.fir 282052:4]
  wire  _T_1 = _io_serial_in_ready_T & io_serial_in_valid; // @[SerialAdapter.scala 138:25 chipyard.TestHarness.RocketConfig.fir 282059:4]
  wire  _GEN_3 = _T_1 ? 1'h0 : idx; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.RocketConfig.fir 282060:4 SerialAdapter.scala 140:9 chipyard.TestHarness.RocketConfig.fir 282062:6 SerialAdapter.scala 91:16 chipyard.TestHarness.RocketConfig.fir 281596:4]
  wire [63:0] _GEN_4 = _T_1 ? 64'h0 : addr; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.RocketConfig.fir 282060:4 SerialAdapter.scala 141:10 chipyard.TestHarness.RocketConfig.fir 282063:6 SerialAdapter.scala 87:17 chipyard.TestHarness.RocketConfig.fir 281592:4]
  wire [63:0] _GEN_5 = _T_1 ? 64'h0 : len; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.RocketConfig.fir 282060:4 SerialAdapter.scala 142:9 chipyard.TestHarness.RocketConfig.fir 282064:6 SerialAdapter.scala 88:16 chipyard.TestHarness.RocketConfig.fir 281593:4]
  wire [3:0] _GEN_6 = _T_1 ? 4'h1 : state; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.RocketConfig.fir 282060:4 SerialAdapter.scala 143:11 chipyard.TestHarness.RocketConfig.fir 282065:6 SerialAdapter.scala 97:22 chipyard.TestHarness.RocketConfig.fir 281597:4]
  wire  _T_3 = _io_serial_in_ready_T_1 & io_serial_in_valid; // @[SerialAdapter.scala 146:26 chipyard.TestHarness.RocketConfig.fir 282068:4]
  wire [5:0] _addr_T = {idx,5'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 282071:6]
  wire [94:0] _GEN_59 = {{63'd0}, io_serial_in_bits}; // @[SerialAdapter.scala 132:12 chipyard.TestHarness.RocketConfig.fir 282072:6]
  wire [94:0] _addr_T_1 = _GEN_59 << _addr_T; // @[SerialAdapter.scala 132:12 chipyard.TestHarness.RocketConfig.fir 282072:6]
  wire [94:0] _GEN_60 = {{31'd0}, addr}; // @[SerialAdapter.scala 147:18 chipyard.TestHarness.RocketConfig.fir 282073:6]
  wire [94:0] _addr_T_2 = _GEN_60 | _addr_T_1; // @[SerialAdapter.scala 147:18 chipyard.TestHarness.RocketConfig.fir 282073:6]
  wire  _idx_T_1 = idx + 1'h1; // @[SerialAdapter.scala 148:16 chipyard.TestHarness.RocketConfig.fir 282076:6]
  wire  _GEN_7 = idx ? 1'h0 : _idx_T_1; // @[SerialAdapter.scala 149:43 chipyard.TestHarness.RocketConfig.fir 282079:6 SerialAdapter.scala 150:11 chipyard.TestHarness.RocketConfig.fir 282080:8 SerialAdapter.scala 148:9 chipyard.TestHarness.RocketConfig.fir 282077:6]
  wire [3:0] _GEN_8 = idx ? 4'h2 : _GEN_6; // @[SerialAdapter.scala 149:43 chipyard.TestHarness.RocketConfig.fir 282079:6 SerialAdapter.scala 151:13 chipyard.TestHarness.RocketConfig.fir 282081:8]
  wire [94:0] _GEN_9 = _T_3 ? _addr_T_2 : {{31'd0}, _GEN_4}; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.RocketConfig.fir 282069:4 SerialAdapter.scala 147:10 chipyard.TestHarness.RocketConfig.fir 282074:6]
  wire  _GEN_10 = _T_3 ? _GEN_7 : _GEN_3; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.RocketConfig.fir 282069:4]
  wire [3:0] _GEN_11 = _T_3 ? _GEN_8 : _GEN_6; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.RocketConfig.fir 282069:4]
  wire  _T_6 = _io_serial_in_ready_T_2 & io_serial_in_valid; // @[SerialAdapter.scala 155:25 chipyard.TestHarness.RocketConfig.fir 282085:4]
  wire [94:0] _GEN_62 = {{31'd0}, len}; // @[SerialAdapter.scala 156:16 chipyard.TestHarness.RocketConfig.fir 282090:6]
  wire [94:0] _len_T_2 = _GEN_62 | _addr_T_1; // @[SerialAdapter.scala 156:16 chipyard.TestHarness.RocketConfig.fir 282090:6]
  wire  _T_8 = cmd == 32'h1; // @[SerialAdapter.scala 160:17 chipyard.TestHarness.RocketConfig.fir 282099:8]
  wire  _T_9 = cmd == 32'h0; // @[SerialAdapter.scala 163:24 chipyard.TestHarness.RocketConfig.fir 282105:10]
  wire  _T_12 = ~reset; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.RocketConfig.fir 282112:12]
  wire [3:0] _GEN_12 = _T_9 ? 4'h3 : _GEN_11; // @[SerialAdapter.scala 163:38 chipyard.TestHarness.RocketConfig.fir 282106:10 SerialAdapter.scala 164:15 chipyard.TestHarness.RocketConfig.fir 282107:12]
  wire [1:0] _GEN_13 = _T_8 ? 2'h0 : bodyValid; // @[SerialAdapter.scala 160:32 chipyard.TestHarness.RocketConfig.fir 282100:8 SerialAdapter.scala 161:19 chipyard.TestHarness.RocketConfig.fir 282101:10 SerialAdapter.scala 90:22 chipyard.TestHarness.RocketConfig.fir 281595:4]
  wire [3:0] _GEN_14 = _T_8 ? 4'h6 : _GEN_12; // @[SerialAdapter.scala 160:32 chipyard.TestHarness.RocketConfig.fir 282100:8 SerialAdapter.scala 162:15 chipyard.TestHarness.RocketConfig.fir 282102:10]
  wire  _GEN_15 = idx ? addr[2] : _idx_T_1; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.RocketConfig.fir 282096:6 SerialAdapter.scala 159:11 chipyard.TestHarness.RocketConfig.fir 282098:8 SerialAdapter.scala 157:9 chipyard.TestHarness.RocketConfig.fir 282094:6]
  wire [1:0] _GEN_16 = idx ? _GEN_13 : bodyValid; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.RocketConfig.fir 282096:6 SerialAdapter.scala 90:22 chipyard.TestHarness.RocketConfig.fir 281595:4]
  wire [3:0] _GEN_17 = idx ? _GEN_14 : _GEN_11; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.RocketConfig.fir 282096:6]
  wire [94:0] _GEN_18 = _T_6 ? _len_T_2 : {{31'd0}, _GEN_5}; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.RocketConfig.fir 282086:4 SerialAdapter.scala 156:9 chipyard.TestHarness.RocketConfig.fir 282091:6]
  wire  _GEN_19 = _T_6 ? _GEN_15 : _GEN_10; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.RocketConfig.fir 282086:4]
  wire [1:0] _GEN_20 = _T_6 ? _GEN_16 : bodyValid; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.RocketConfig.fir 282086:4 SerialAdapter.scala 90:22 chipyard.TestHarness.RocketConfig.fir 281595:4]
  wire [3:0] _GEN_21 = _T_6 ? _GEN_17 : _GEN_11; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.RocketConfig.fir 282086:4]
  wire  _T_14 = _bundleOut_0_a_valid_T_1 & auto_out_a_ready; // @[SerialAdapter.scala 171:30 chipyard.TestHarness.RocketConfig.fir 282121:4]
  wire [3:0] _GEN_22 = _T_14 ? 4'h4 : _GEN_21; // @[SerialAdapter.scala 171:46 chipyard.TestHarness.RocketConfig.fir 282122:4 SerialAdapter.scala 172:11 chipyard.TestHarness.RocketConfig.fir 282123:6]
  wire  _T_16 = _bundleOut_0_d_ready_T_1 & auto_out_d_valid; // @[SerialAdapter.scala 175:31 chipyard.TestHarness.RocketConfig.fir 282126:4]
  wire [31:0] _GEN_23 = _T_16 ? auto_out_d_bits_data[31:0] : body_0; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.RocketConfig.fir 282127:4 SerialAdapter.scala 176:10 chipyard.TestHarness.RocketConfig.fir 282135:6 SerialAdapter.scala 89:17 chipyard.TestHarness.RocketConfig.fir 281594:4]
  wire [31:0] _GEN_24 = _T_16 ? auto_out_d_bits_data[63:32] : body_1; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.RocketConfig.fir 282127:4 SerialAdapter.scala 176:10 chipyard.TestHarness.RocketConfig.fir 282136:6 SerialAdapter.scala 89:17 chipyard.TestHarness.RocketConfig.fir 281594:4]
  wire  _GEN_25 = _T_16 ? addr[2] : _GEN_19; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.RocketConfig.fir 282127:4 SerialAdapter.scala 177:9 chipyard.TestHarness.RocketConfig.fir 282138:6]
  wire [94:0] _GEN_26 = _T_16 ? {{63'd0}, nextAddr} : _GEN_9; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.RocketConfig.fir 282127:4 SerialAdapter.scala 178:10 chipyard.TestHarness.RocketConfig.fir 282139:6]
  wire [3:0] _GEN_27 = _T_16 ? 4'h5 : _GEN_22; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.RocketConfig.fir 282127:4 SerialAdapter.scala 179:11 chipyard.TestHarness.RocketConfig.fir 282140:6]
  wire  _T_20 = _io_serial_out_valid_T & io_serial_out_ready; // @[SerialAdapter.scala 182:31 chipyard.TestHarness.RocketConfig.fir 282143:4]
  wire [63:0] _len_T_4 = len - 64'h1; // @[SerialAdapter.scala 184:16 chipyard.TestHarness.RocketConfig.fir 282149:6]
  wire  _T_21 = len == 64'h0; // @[SerialAdapter.scala 185:15 chipyard.TestHarness.RocketConfig.fir 282151:6]
  wire [3:0] _GEN_28 = idx ? 4'h3 : _GEN_27; // @[SerialAdapter.scala 186:48 chipyard.TestHarness.RocketConfig.fir 282157:8 SerialAdapter.scala 186:56 chipyard.TestHarness.RocketConfig.fir 282158:10]
  wire [3:0] _GEN_29 = _T_21 ? 4'h0 : _GEN_28; // @[SerialAdapter.scala 185:24 chipyard.TestHarness.RocketConfig.fir 282152:6 SerialAdapter.scala 185:32 chipyard.TestHarness.RocketConfig.fir 282153:8]
  wire  _GEN_30 = _T_20 ? _idx_T_1 : _GEN_25; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.RocketConfig.fir 282144:4 SerialAdapter.scala 183:9 chipyard.TestHarness.RocketConfig.fir 282147:6]
  wire [94:0] _GEN_31 = _T_20 ? {{31'd0}, _len_T_4} : _GEN_18; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.RocketConfig.fir 282144:4 SerialAdapter.scala 184:9 chipyard.TestHarness.RocketConfig.fir 282150:6]
  wire [3:0] _GEN_32 = _T_20 ? _GEN_29 : _GEN_27; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.RocketConfig.fir 282144:4]
  wire  _T_24 = _io_serial_in_ready_T_3 & io_serial_in_valid; // @[SerialAdapter.scala 189:32 chipyard.TestHarness.RocketConfig.fir 282162:4]
  wire [1:0] _bodyValid_T = 2'h1 << idx; // @[OneHot.scala 58:35 chipyard.TestHarness.RocketConfig.fir 282165:6]
  wire [1:0] _bodyValid_T_1 = bodyValid | _bodyValid_T; // @[SerialAdapter.scala 191:28 chipyard.TestHarness.RocketConfig.fir 282166:6]
  wire  _T_27 = idx | _T_21; // @[SerialAdapter.scala 192:42 chipyard.TestHarness.RocketConfig.fir 282170:6]
  wire [3:0] _GEN_35 = _T_27 ? 4'h7 : _GEN_32; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.RocketConfig.fir 282171:6 SerialAdapter.scala 193:13 chipyard.TestHarness.RocketConfig.fir 282172:8]
  wire  _GEN_36 = _T_27 ? _GEN_30 : _idx_T_1; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.RocketConfig.fir 282171:6 SerialAdapter.scala 195:11 chipyard.TestHarness.RocketConfig.fir 282177:8]
  wire [94:0] _GEN_37 = _T_27 ? _GEN_31 : {{31'd0}, _len_T_4}; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.RocketConfig.fir 282171:6 SerialAdapter.scala 196:11 chipyard.TestHarness.RocketConfig.fir 282180:8]
  wire [1:0] _GEN_40 = _T_24 ? _bodyValid_T_1 : _GEN_20; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.RocketConfig.fir 282163:4 SerialAdapter.scala 191:15 chipyard.TestHarness.RocketConfig.fir 282167:6]
  wire  _GEN_42 = _T_24 ? _GEN_36 : _GEN_30; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.RocketConfig.fir 282163:4]
  wire [94:0] _GEN_43 = _T_24 ? _GEN_37 : _GEN_31; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.RocketConfig.fir 282163:4]
  wire  _T_29 = _bundleOut_0_a_valid_T & auto_out_a_ready; // @[SerialAdapter.scala 200:32 chipyard.TestHarness.RocketConfig.fir 282184:4]
  wire  _T_31 = _bundleOut_0_d_ready_T & auto_out_d_valid; // @[SerialAdapter.scala 204:31 chipyard.TestHarness.RocketConfig.fir 282189:4]
  wire [94:0] _GEN_46 = _T_21 ? _GEN_26 : {{63'd0}, nextAddr}; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.RocketConfig.fir 282192:6 SerialAdapter.scala 208:12 chipyard.TestHarness.RocketConfig.fir 282196:8]
  wire [94:0] _GEN_47 = _T_21 ? _GEN_43 : {{31'd0}, _len_T_4}; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.RocketConfig.fir 282192:6 SerialAdapter.scala 209:11 chipyard.TestHarness.RocketConfig.fir 282199:8]
  wire  _GEN_48 = _T_21 & _GEN_42; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.RocketConfig.fir 282192:6 SerialAdapter.scala 210:11 chipyard.TestHarness.RocketConfig.fir 282200:8]
  wire [94:0] _GEN_51 = _T_31 ? _GEN_46 : _GEN_26; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.RocketConfig.fir 282190:4]
  wire [94:0] _GEN_52 = _T_31 ? _GEN_47 : _GEN_43; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.RocketConfig.fir 282190:4]
  wire  _GEN_67 = _T_6 & idx & ~_T_8 & ~_T_9; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.RocketConfig.fir 282114:14]
  assign auto_out_a_valid = _bundleOut_0_a_valid_T | _bundleOut_0_a_valid_T_1; // @[package.scala 72:59 chipyard.TestHarness.RocketConfig.fir 282033:4]
  assign auto_out_a_bits_opcode = _bundleOut_0_a_valid_T ? 3'h1 : 3'h4; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.RocketConfig.fir 282036:4]
  assign auto_out_a_bits_size = _bundleOut_0_a_valid_T ? 4'h3 : get_acquire_size; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.RocketConfig.fir 282036:4]
  assign auto_out_a_bits_address = _bundleOut_0_a_valid_T ? put_acquire_address : get_acquire_address; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.RocketConfig.fir 282036:4]
  assign auto_out_a_bits_mask = _bundleOut_0_a_valid_T ? wmask : get_acquire_mask; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.RocketConfig.fir 282036:4]
  assign auto_out_a_bits_data = _bundleOut_0_a_valid_T ? put_acquire_data : 64'h0; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.RocketConfig.fir 282036:4]
  assign auto_out_d_ready = _bundleOut_0_d_ready_T | _bundleOut_0_d_ready_T_1; // @[package.scala 72:59 chipyard.TestHarness.RocketConfig.fir 282053:4]
  assign io_serial_in_ready = _io_serial_in_ready_T_5 | _io_serial_in_ready_T_3; // @[package.scala 72:59 chipyard.TestHarness.RocketConfig.fir 281604:4]
  assign io_serial_out_valid = state == 4'h5; // @[SerialAdapter.scala 100:32 chipyard.TestHarness.RocketConfig.fir 281606:4]
  assign io_serial_out_bits = idx ? body_1 : body_0; // @[SerialAdapter.scala 101:22 chipyard.TestHarness.RocketConfig.fir 281608:4 SerialAdapter.scala 101:22 chipyard.TestHarness.RocketConfig.fir 281608:4]
  always @(posedge clock) begin
    if (_T_1) begin // @[SerialAdapter.scala 138:48 chipyard.TestHarness.RocketConfig.fir 282060:4]
      cmd <= io_serial_in_bits; // @[SerialAdapter.scala 139:9 chipyard.TestHarness.RocketConfig.fir 282061:6]
    end
    addr <= _GEN_51[63:0];
    len <= _GEN_52[63:0];
    if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.RocketConfig.fir 282163:4]
      if (~idx) begin // @[SerialAdapter.scala 190:15 chipyard.TestHarness.RocketConfig.fir 282164:6]
        body_0 <= io_serial_in_bits; // @[SerialAdapter.scala 190:15 chipyard.TestHarness.RocketConfig.fir 282164:6]
      end else begin
        body_0 <= _GEN_23;
      end
    end else begin
      body_0 <= _GEN_23;
    end
    if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.RocketConfig.fir 282163:4]
      if (idx) begin // @[SerialAdapter.scala 190:15 chipyard.TestHarness.RocketConfig.fir 282164:6]
        body_1 <= io_serial_in_bits; // @[SerialAdapter.scala 190:15 chipyard.TestHarness.RocketConfig.fir 282164:6]
      end else begin
        body_1 <= _GEN_24;
      end
    end else begin
      body_1 <= _GEN_24;
    end
    if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.RocketConfig.fir 282190:4]
      if (_T_21) begin // @[SerialAdapter.scala 205:24 chipyard.TestHarness.RocketConfig.fir 282192:6]
        bodyValid <= _GEN_40;
      end else begin
        bodyValid <= 2'h0; // @[SerialAdapter.scala 211:17 chipyard.TestHarness.RocketConfig.fir 282201:8]
      end
    end else begin
      bodyValid <= _GEN_40;
    end
    if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.RocketConfig.fir 282190:4]
      idx <= _GEN_48;
    end else if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.RocketConfig.fir 282163:4]
      if (_T_27) begin // @[SerialAdapter.scala 192:58 chipyard.TestHarness.RocketConfig.fir 282171:6]
        idx <= _GEN_30;
      end else begin
        idx <= _idx_T_1; // @[SerialAdapter.scala 195:11 chipyard.TestHarness.RocketConfig.fir 282177:8]
      end
    end else begin
      idx <= _GEN_30;
    end
    if (reset) begin // @[SerialAdapter.scala 97:22 chipyard.TestHarness.RocketConfig.fir 281597:4]
      state <= 4'h0; // @[SerialAdapter.scala 97:22 chipyard.TestHarness.RocketConfig.fir 281597:4]
    end else if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.RocketConfig.fir 282190:4]
      if (_T_21) begin // @[SerialAdapter.scala 205:24 chipyard.TestHarness.RocketConfig.fir 282192:6]
        state <= 4'h0; // @[SerialAdapter.scala 206:13 chipyard.TestHarness.RocketConfig.fir 282193:8]
      end else begin
        state <= 4'h6; // @[SerialAdapter.scala 212:13 chipyard.TestHarness.RocketConfig.fir 282202:8]
      end
    end else if (_T_29) begin // @[SerialAdapter.scala 200:48 chipyard.TestHarness.RocketConfig.fir 282185:4]
      state <= 4'h8; // @[SerialAdapter.scala 201:11 chipyard.TestHarness.RocketConfig.fir 282186:6]
    end else if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.RocketConfig.fir 282163:4]
      state <= _GEN_35;
    end else begin
      state <= _GEN_32;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & idx & ~_T_8 & ~_T_9 & _T_12) begin
          $fwrite(32'h80000002,
            "Assertion failed: Bad TSI command\n    at SerialAdapter.scala:166 assert(false.B, \"Bad TSI command\")\n"); // @[SerialAdapter.scala 166:15 chipyard.TestHarness.RocketConfig.fir 282114:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_12) begin
          $fatal; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.RocketConfig.fir 282115:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cmd = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  addr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  len = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  body_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  body_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bodyValid = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  idx = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_53_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 282222:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 282223:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 282224:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input  [3:0]  io_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input         io_in_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input  [31:0] io_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input  [3:0]  io_in_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input         io_in_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input  [2:0]  io_in_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 282225:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 284164:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 284471:4]
  wire  _source_ok_T = ~io_in_a_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.RocketConfig.fir 282236:6]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 282241:6]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 282243:6]
  wire [31:0] _GEN_71 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.RocketConfig.fir 282244:6]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.RocketConfig.fir 282244:6]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24 chipyard.TestHarness.RocketConfig.fir 282245:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.RocketConfig.fir 282247:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.RocketConfig.fir 282248:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.RocketConfig.fir 282250:6]
  wire  _mask_T = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21 chipyard.TestHarness.RocketConfig.fir 282251:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 282252:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 282253:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 282254:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282256:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282257:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282259:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282260:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 282261:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 282262:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 282263:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282264:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282265:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282266:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282267:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282268:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282269:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282270:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282271:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282272:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282273:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282274:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282275:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 282276:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 282277:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 282278:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282279:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282280:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282281:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282282:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282283:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282284:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282285:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282286:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282287:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282288:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282289:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282290:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282291:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282292:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282293:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282294:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282295:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282296:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282297:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282298:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282299:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 282300:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 282301:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 282302:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 282309:6]
  wire [32:0] _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 282313:6]
  wire  _T_15 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.RocketConfig.fir 282325:6]
  wire  _T_17 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42 chipyard.TestHarness.RocketConfig.fir 282328:8]
  wire  _T_20 = _T_17 & _source_ok_T; // @[Parameters.scala 1160:30 chipyard.TestHarness.RocketConfig.fir 282331:8]
  wire [32:0] _T_26 = $signed(_T_7) & -33'sh101000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 282337:8]
  wire  _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 282338:8]
  wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 282339:8]
  wire [32:0] _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 282340:8]
  wire [32:0] _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 282342:8]
  wire  _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 282343:8]
  wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 282344:8]
  wire [32:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 282345:8]
  wire [32:0] _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 282347:8]
  wire  _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 282348:8]
  wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 282349:8]
  wire [32:0] _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 282350:8]
  wire [32:0] _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 282352:8]
  wire  _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 282353:8]
  wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h2010000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 282354:8]
  wire [32:0] _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 282355:8]
  wire [32:0] _T_46 = $signed(_T_44) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 282357:8]
  wire  _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 282358:8]
  wire [31:0] _T_48 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 282359:8]
  wire [32:0] _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 282360:8]
  wire [32:0] _T_51 = $signed(_T_49) & -33'sh4000000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 282362:8]
  wire  _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 282363:8]
  wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h54000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 282364:8]
  wire [32:0] _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 282365:8]
  wire [32:0] _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 282367:8]
  wire  _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 282368:8]
  wire  _T_58 = _T_27 | _T_32; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282369:8]
  wire  _T_65 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48 chipyard.TestHarness.RocketConfig.fir 282376:8]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 282378:8]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 282379:8]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 282381:8]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 282382:8]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 282383:8]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 282384:8]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh10000000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 282386:8]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 282387:8]
  wire  _T_77 = _T_71 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282388:8]
  wire  _T_78 = _T_65 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 282389:8]
  wire  _T_81 = _T_20 & _T_78; // @[Monitor.scala 82:72 chipyard.TestHarness.RocketConfig.fir 282392:8]
  wire  _T_83 = _T_81 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282394:8]
  wire  _T_84 = ~_T_83; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282395:8]
  wire  _T_147 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282462:8]
  wire  _T_149 = _source_ok_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282468:8]
  wire  _T_150 = ~_T_149; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282469:8]
  wire  _T_153 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282476:8]
  wire  _T_154 = ~_T_153; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282477:8]
  wire  _T_156 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282483:8]
  wire  _T_157 = ~_T_156; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282484:8]
  wire  _T_158 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.RocketConfig.fir 282489:8]
  wire  _T_160 = _T_158 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282491:8]
  wire  _T_161 = ~_T_160; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282492:8]
  wire [7:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.RocketConfig.fir 282497:8]
  wire  _T_163 = _T_162 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.RocketConfig.fir 282498:8]
  wire  _T_165 = _T_163 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282500:8]
  wire  _T_166 = ~_T_165; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282501:8]
  wire  _T_167 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.RocketConfig.fir 282506:8]
  wire  _T_169 = _T_167 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282508:8]
  wire  _T_170 = ~_T_169; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282509:8]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.RocketConfig.fir 282515:6]
  wire  _T_318 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.RocketConfig.fir 282687:8]
  wire  _T_320 = _T_318 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282689:8]
  wire  _T_321 = ~_T_320; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282690:8]
  wire  _T_331 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.RocketConfig.fir 282713:6]
  wire  _T_339 = _T_20 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282722:8]
  wire  _T_340 = ~_T_339; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282723:8]
  wire  _T_350 = _T_17 & _T_32; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 282737:8]
  wire  _T_352 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.RocketConfig.fir 282739:8]
  wire  _T_395 = _T_27 | _T_37; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282782:8]
  wire  _T_396 = _T_395 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282783:8]
  wire  _T_397 = _T_396 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282784:8]
  wire  _T_398 = _T_397 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282785:8]
  wire  _T_399 = _T_398 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282786:8]
  wire  _T_400 = _T_399 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282787:8]
  wire  _T_401 = _T_400 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282788:8]
  wire  _T_402 = _T_352 & _T_401; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 282789:8]
  wire  _T_404 = _T_350 | _T_402; // @[Parameters.scala 672:30 chipyard.TestHarness.RocketConfig.fir 282791:8]
  wire  _T_406 = _T_404 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282793:8]
  wire  _T_407 = ~_T_406; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282794:8]
  wire  _T_414 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.RocketConfig.fir 282813:8]
  wire  _T_416 = _T_414 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282815:8]
  wire  _T_417 = ~_T_416; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282816:8]
  wire  _T_418 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.RocketConfig.fir 282821:8]
  wire  _T_420 = _T_418 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282823:8]
  wire  _T_421 = ~_T_420; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282824:8]
  wire  _T_426 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.RocketConfig.fir 282838:6]
  wire  _T_482 = _T_27 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282895:8]
  wire  _T_483 = _T_482 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282896:8]
  wire  _T_484 = _T_483 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282897:8]
  wire  _T_485 = _T_484 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282898:8]
  wire  _T_486 = _T_485 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282899:8]
  wire  _T_487 = _T_486 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 282900:8]
  wire  _T_488 = _T_352 & _T_487; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 282901:8]
  wire  _T_497 = _T_350 | _T_488; // @[Parameters.scala 672:30 chipyard.TestHarness.RocketConfig.fir 282910:8]
  wire  _T_499 = _T_20 & _T_497; // @[Monitor.scala 115:71 chipyard.TestHarness.RocketConfig.fir 282912:8]
  wire  _T_501 = _T_499 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282914:8]
  wire  _T_502 = ~_T_501; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282915:8]
  wire  _T_517 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.RocketConfig.fir 282951:6]
  wire [7:0] _T_604 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.RocketConfig.fir 283055:8]
  wire [7:0] _T_605 = io_in_a_bits_mask & _T_604; // @[Monitor.scala 127:31 chipyard.TestHarness.RocketConfig.fir 283056:8]
  wire  _T_606 = _T_605 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.RocketConfig.fir 283057:8]
  wire  _T_608 = _T_606 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283059:8]
  wire  _T_609 = ~_T_608; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283060:8]
  wire  _T_610 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.RocketConfig.fir 283066:6]
  wire  _T_618 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 92:42 chipyard.TestHarness.RocketConfig.fir 283075:8]
  wire  _T_662 = _T_58 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 283119:8]
  wire  _T_663 = _T_662 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 283120:8]
  wire  _T_664 = _T_663 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 283121:8]
  wire  _T_665 = _T_664 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 283122:8]
  wire  _T_666 = _T_665 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 283123:8]
  wire  _T_667 = _T_666 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 283124:8]
  wire  _T_668 = _T_618 & _T_667; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 283125:8]
  wire  _T_678 = _T_20 & _T_668; // @[Monitor.scala 131:74 chipyard.TestHarness.RocketConfig.fir 283135:8]
  wire  _T_680 = _T_678 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283137:8]
  wire  _T_681 = ~_T_680; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283138:8]
  wire  _T_688 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.RocketConfig.fir 283157:8]
  wire  _T_690 = _T_688 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283159:8]
  wire  _T_691 = ~_T_690; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283160:8]
  wire  _T_696 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.RocketConfig.fir 283174:6]
  wire  _T_774 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.RocketConfig.fir 283265:8]
  wire  _T_776 = _T_774 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283267:8]
  wire  _T_777 = ~_T_776; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283268:8]
  wire  _T_782 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.RocketConfig.fir 283282:6]
  wire  _T_851 = _T_352 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 283352:8]
  wire  _T_854 = _T_350 | _T_851; // @[Parameters.scala 672:30 chipyard.TestHarness.RocketConfig.fir 283355:8]
  wire  _T_855 = _T_20 & _T_854; // @[Monitor.scala 147:68 chipyard.TestHarness.RocketConfig.fir 283356:8]
  wire  _T_857 = _T_855 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283358:8]
  wire  _T_858 = ~_T_857; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283359:8]
  wire  _T_865 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.RocketConfig.fir 283378:8]
  wire  _T_867 = _T_865 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283380:8]
  wire  _T_868 = ~_T_867; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283381:8]
  wire  _T_877 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.RocketConfig.fir 283405:6]
  wire  _T_879 = _T_877 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283407:6]
  wire  _T_880 = ~_T_879; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283408:6]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.RocketConfig.fir 283413:6]
  wire  _T_881 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.RocketConfig.fir 283418:6]
  wire  _T_883 = _source_ok_T_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283421:8]
  wire  _T_884 = ~_T_883; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283422:8]
  wire  _T_885 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.RocketConfig.fir 283427:8]
  wire  _T_887 = _T_885 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283429:8]
  wire  _T_888 = ~_T_887; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283430:8]
  wire  _T_889 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.RocketConfig.fir 283435:8]
  wire  _T_891 = _T_889 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283437:8]
  wire  _T_892 = ~_T_891; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283438:8]
  wire  _T_893 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.RocketConfig.fir 283443:8]
  wire  _T_895 = _T_893 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283445:8]
  wire  _T_896 = ~_T_895; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283446:8]
  wire  _T_897 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.RocketConfig.fir 283451:8]
  wire  _T_899 = _T_897 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283453:8]
  wire  _T_900 = ~_T_899; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283454:8]
  wire  _T_901 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.RocketConfig.fir 283460:6]
  wire  _T_912 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.RocketConfig.fir 283484:8]
  wire  _T_914 = _T_912 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283486:8]
  wire  _T_915 = ~_T_914; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283487:8]
  wire  _T_916 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.RocketConfig.fir 283492:8]
  wire  _T_918 = _T_916 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283494:8]
  wire  _T_919 = ~_T_918; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283495:8]
  wire  _T_929 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.RocketConfig.fir 283518:6]
  wire  _T_949 = _T_897 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.RocketConfig.fir 283559:8]
  wire  _T_951 = _T_949 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283561:8]
  wire  _T_952 = ~_T_951; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283562:8]
  wire  _T_958 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.RocketConfig.fir 283577:6]
  wire  _T_975 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.RocketConfig.fir 283612:6]
  wire  _T_993 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.RocketConfig.fir 283648:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 283714:4]
  wire [8:0] a_first_beats1_decode = is_aligned_mask[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.RocketConfig.fir 283719:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.RocketConfig.fir 283721:4]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283723:4]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 283725:4]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 283726:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.RocketConfig.fir 283737:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.RocketConfig.fir 283738:4]
  reg [3:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.RocketConfig.fir 283739:4]
  reg  source; // @[Monitor.scala 387:22 chipyard.TestHarness.RocketConfig.fir 283740:4]
  reg [31:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.RocketConfig.fir 283741:4]
  wire  _T_1022 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.RocketConfig.fir 283742:4]
  wire  _T_1023 = io_in_a_valid & _T_1022; // @[Monitor.scala 389:19 chipyard.TestHarness.RocketConfig.fir 283743:4]
  wire  _T_1024 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.RocketConfig.fir 283745:6]
  wire  _T_1026 = _T_1024 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283747:6]
  wire  _T_1027 = ~_T_1026; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283748:6]
  wire  _T_1028 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.RocketConfig.fir 283753:6]
  wire  _T_1030 = _T_1028 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283755:6]
  wire  _T_1031 = ~_T_1030; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283756:6]
  wire  _T_1032 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.RocketConfig.fir 283761:6]
  wire  _T_1034 = _T_1032 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283763:6]
  wire  _T_1035 = ~_T_1034; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283764:6]
  wire  _T_1036 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.RocketConfig.fir 283769:6]
  wire  _T_1038 = _T_1036 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283771:6]
  wire  _T_1039 = ~_T_1038; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283772:6]
  wire  _T_1040 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.RocketConfig.fir 283777:6]
  wire  _T_1042 = _T_1040 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283779:6]
  wire  _T_1043 = ~_T_1042; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283780:6]
  wire  _T_1045 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.RocketConfig.fir 283787:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 283795:4]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 283797:4]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 283799:4]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.RocketConfig.fir 283800:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.RocketConfig.fir 283801:4]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283803:4]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 283805:4]
  wire  d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 283806:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.RocketConfig.fir 283817:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.RocketConfig.fir 283818:4]
  reg [3:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.RocketConfig.fir 283819:4]
  reg  source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.RocketConfig.fir 283820:4]
  reg [2:0] sink; // @[Monitor.scala 539:22 chipyard.TestHarness.RocketConfig.fir 283821:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.RocketConfig.fir 283822:4]
  wire  _T_1046 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.RocketConfig.fir 283823:4]
  wire  _T_1047 = io_in_d_valid & _T_1046; // @[Monitor.scala 541:19 chipyard.TestHarness.RocketConfig.fir 283824:4]
  wire  _T_1048 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.RocketConfig.fir 283826:6]
  wire  _T_1050 = _T_1048 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283828:6]
  wire  _T_1051 = ~_T_1050; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283829:6]
  wire  _T_1052 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.RocketConfig.fir 283834:6]
  wire  _T_1054 = _T_1052 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283836:6]
  wire  _T_1055 = ~_T_1054; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283837:6]
  wire  _T_1056 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.RocketConfig.fir 283842:6]
  wire  _T_1058 = _T_1056 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283844:6]
  wire  _T_1059 = ~_T_1058; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283845:6]
  wire  _T_1060 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.RocketConfig.fir 283850:6]
  wire  _T_1062 = _T_1060 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283852:6]
  wire  _T_1063 = ~_T_1062; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283853:6]
  wire  _T_1064 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.RocketConfig.fir 283858:6]
  wire  _T_1066 = _T_1064 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283860:6]
  wire  _T_1067 = ~_T_1066; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283861:6]
  wire  _T_1068 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.RocketConfig.fir 283866:6]
  wire  _T_1070 = _T_1068 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283868:6]
  wire  _T_1071 = ~_T_1070; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283869:6]
  wire  _T_1073 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.RocketConfig.fir 283876:4]
  reg  inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 283885:4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 283886:4]
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 283887:4]
  reg [8:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283897:4]
  wire [8:0] a_first_counter1_1 = a_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 283899:4]
  wire  a_first_1 = a_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 283900:4]
  reg [8:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283919:4]
  wire [8:0] d_first_counter1_1 = d_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 283921:4]
  wire  d_first_1 = d_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 283922:4]
  wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.RocketConfig.fir 283943:4]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.RocketConfig.fir 283943:4]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.RocketConfig.fir 283944:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.RocketConfig.fir 283948:4]
  wire [15:0] _GEN_73 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.RocketConfig.fir 283949:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.RocketConfig.fir 283949:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.RocketConfig.fir 283950:4]
  wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65 chipyard.TestHarness.RocketConfig.fir 283954:4]
  wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.RocketConfig.fir 283955:4]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.RocketConfig.fir 283959:4]
  wire [15:0] _GEN_75 = {{8'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.RocketConfig.fir 283960:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.RocketConfig.fir 283960:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.RocketConfig.fir 283961:4]
  wire  _T_1074 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.RocketConfig.fir 283985:4]
  wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.RocketConfig.fir 283988:6]
  wire [1:0] _GEN_15 = _T_1074 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.RocketConfig.fir 283987:4 Monitor.scala 649:22 chipyard.TestHarness.RocketConfig.fir 283989:6 chipyard.TestHarness.RocketConfig.fir 283936:4]
  wire  _T_1077 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.RocketConfig.fir 283992:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.RocketConfig.fir 283997:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.RocketConfig.fir 283998:6]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.RocketConfig.fir 284000:6]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.RocketConfig.fir 284001:6]
  wire [2:0] _GEN_77 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.RocketConfig.fir 284003:6]
  wire [3:0] _a_opcodes_set_T = {{1'd0}, _GEN_77}; // @[Monitor.scala 656:79 chipyard.TestHarness.RocketConfig.fir 284003:6]
  wire [3:0] a_opcodes_set_interm = _T_1077 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 283994:4 Monitor.scala 654:28 chipyard.TestHarness.RocketConfig.fir 283999:6 chipyard.TestHarness.RocketConfig.fir 283982:4]
  wire [18:0] _GEN_78 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.RocketConfig.fir 284004:6]
  wire [18:0] _a_opcodes_set_T_1 = _GEN_78 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.RocketConfig.fir 284004:6]
  wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 657:77 chipyard.TestHarness.RocketConfig.fir 284006:6]
  wire [4:0] a_sizes_set_interm = _T_1077 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 283994:4 Monitor.scala 655:28 chipyard.TestHarness.RocketConfig.fir 284002:6 chipyard.TestHarness.RocketConfig.fir 283984:4]
  wire [19:0] _GEN_79 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.RocketConfig.fir 284007:6]
  wire [19:0] _a_sizes_set_T_1 = _GEN_79 << _a_sizes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.RocketConfig.fir 284007:6]
  wire  _T_1079 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.RocketConfig.fir 284009:6]
  wire  _T_1081 = ~_T_1079; // @[Monitor.scala 658:17 chipyard.TestHarness.RocketConfig.fir 284011:6]
  wire  _T_1083 = _T_1081 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 284013:6]
  wire  _T_1084 = ~_T_1083; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 284014:6]
  wire [1:0] _GEN_16 = _T_1077 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 283994:4 Monitor.scala 653:28 chipyard.TestHarness.RocketConfig.fir 283996:6 chipyard.TestHarness.RocketConfig.fir 283934:4]
  wire [18:0] _GEN_19 = _T_1077 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 283994:4 Monitor.scala 656:28 chipyard.TestHarness.RocketConfig.fir 284005:6 chipyard.TestHarness.RocketConfig.fir 283938:4]
  wire [19:0] _GEN_20 = _T_1077 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 283994:4 Monitor.scala 657:28 chipyard.TestHarness.RocketConfig.fir 284008:6 chipyard.TestHarness.RocketConfig.fir 283940:4]
  wire  _T_1085 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.RocketConfig.fir 284029:4]
  wire  _T_1087 = ~_T_881; // @[Monitor.scala 671:74 chipyard.TestHarness.RocketConfig.fir 284031:4]
  wire  _T_1088 = _T_1085 & _T_1087; // @[Monitor.scala 671:71 chipyard.TestHarness.RocketConfig.fir 284032:4]
  wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.RocketConfig.fir 284034:6]
  wire [1:0] _GEN_21 = _T_1088 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.RocketConfig.fir 284033:4 Monitor.scala 672:22 chipyard.TestHarness.RocketConfig.fir 284035:6 chipyard.TestHarness.RocketConfig.fir 284023:4]
  wire  _T_1090 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.RocketConfig.fir 284038:4]
  wire  _T_1093 = _T_1090 & _T_1087; // @[Monitor.scala 675:72 chipyard.TestHarness.RocketConfig.fir 284041:4]
  wire [30:0] _GEN_81 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.RocketConfig.fir 284050:6]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_81 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.RocketConfig.fir 284050:6]
  wire [30:0] _GEN_82 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74 chipyard.TestHarness.RocketConfig.fir 284057:6]
  wire [30:0] _d_sizes_clr_T_5 = _GEN_82 << _a_size_lookup_T; // @[Monitor.scala 678:74 chipyard.TestHarness.RocketConfig.fir 284057:6]
  wire [1:0] _GEN_22 = _T_1093 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 284042:4 Monitor.scala 676:21 chipyard.TestHarness.RocketConfig.fir 284044:6 chipyard.TestHarness.RocketConfig.fir 284021:4]
  wire [30:0] _GEN_23 = _T_1093 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 284042:4 Monitor.scala 677:21 chipyard.TestHarness.RocketConfig.fir 284051:6 chipyard.TestHarness.RocketConfig.fir 284025:4]
  wire [30:0] _GEN_24 = _T_1093 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 284042:4 Monitor.scala 678:21 chipyard.TestHarness.RocketConfig.fir 284058:6 chipyard.TestHarness.RocketConfig.fir 284027:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.RocketConfig.fir 284067:6]
  wire  same_cycle_resp = _T_1074 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.RocketConfig.fir 284068:6]
  wire  _T_1098 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.RocketConfig.fir 284069:6]
  wire  _T_1100 = _T_1098 | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.RocketConfig.fir 284071:6]
  wire  _T_1102 = _T_1100 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284073:6]
  wire  _T_1103 = ~_T_1102; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284074:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8]
  wire  _T_1104 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 284080:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 284081:8 Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 284081:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 284081:8 Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 284081:8]
  wire  _T_1105 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 284081:8]
  wire  _T_1106 = _T_1104 | _T_1105; // @[Monitor.scala 685:77 chipyard.TestHarness.RocketConfig.fir 284082:8]
  wire  _T_1108 = _T_1106 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284084:8]
  wire  _T_1109 = ~_T_1108; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284085:8]
  wire  _T_1110 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.RocketConfig.fir 284090:8]
  wire  _T_1112 = _T_1110 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284092:8]
  wire  _T_1113 = ~_T_1112; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284093:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 283941:4 Monitor.scala 634:21 chipyard.TestHarness.RocketConfig.fir 283951:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8]
  wire  _T_1115 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 284101:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 284103:8 Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 284103:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 284103:8 Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 284103:8]
  wire  _T_1117 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 284103:8]
  wire  _T_1118 = _T_1115 | _T_1117; // @[Monitor.scala 689:72 chipyard.TestHarness.RocketConfig.fir 284104:8]
  wire  _T_1120 = _T_1118 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284106:8]
  wire  _T_1121 = ~_T_1120; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284107:8]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.RocketConfig.fir 283952:4 Monitor.scala 638:19 chipyard.TestHarness.RocketConfig.fir 283962:4]
  wire [7:0] _GEN_83 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.RocketConfig.fir 284112:8]
  wire  _T_1122 = _GEN_83 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.RocketConfig.fir 284112:8]
  wire  _T_1124 = _T_1122 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284114:8]
  wire  _T_1125 = ~_T_1124; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284115:8]
  wire  _T_1127 = _T_1085 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.RocketConfig.fir 284123:4]
  wire  _T_1128 = _T_1127 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.RocketConfig.fir 284124:4]
  wire  _T_1130 = _T_1128 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.RocketConfig.fir 284126:4]
  wire  _T_1132 = _T_1130 & _T_1087; // @[Monitor.scala 694:116 chipyard.TestHarness.RocketConfig.fir 284128:4]
  wire  _T_1133 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.RocketConfig.fir 284130:6]
  wire  _T_1134 = _T_1133 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.RocketConfig.fir 284131:6]
  wire  _T_1136 = _T_1134 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284133:6]
  wire  _T_1137 = ~_T_1136; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284134:6]
  wire  a_set_wo_ready = _GEN_15[0]; // @[chipyard.TestHarness.RocketConfig.fir 283935:4]
  wire  d_clr_wo_ready = _GEN_21[0]; // @[chipyard.TestHarness.RocketConfig.fir 284022:4]
  wire  _T_1138 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.RocketConfig.fir 284140:4]
  wire  _T_1139 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.RocketConfig.fir 284141:4]
  wire  _T_1140 = ~_T_1139; // @[Monitor.scala 699:51 chipyard.TestHarness.RocketConfig.fir 284142:4]
  wire  _T_1141 = _T_1138 | _T_1140; // @[Monitor.scala 699:48 chipyard.TestHarness.RocketConfig.fir 284143:4]
  wire  _T_1143 = _T_1141 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284145:4]
  wire  _T_1144 = ~_T_1143; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284146:4]
  wire  a_set = _GEN_16[0]; // @[chipyard.TestHarness.RocketConfig.fir 283933:4]
  wire  _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.RocketConfig.fir 284151:4]
  wire  d_clr = _GEN_22[0]; // @[chipyard.TestHarness.RocketConfig.fir 284020:4]
  wire  _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.RocketConfig.fir 284152:4]
  wire  _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.RocketConfig.fir 284153:4]
  wire [3:0] a_opcodes_set = _GEN_19[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 283937:4]
  wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.RocketConfig.fir 284155:4]
  wire [3:0] d_opcodes_clr = _GEN_23[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 284024:4]
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.RocketConfig.fir 284156:4]
  wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.RocketConfig.fir 284157:4]
  wire [7:0] a_sizes_set = _GEN_20[7:0]; // @[chipyard.TestHarness.RocketConfig.fir 283939:4]
  wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.RocketConfig.fir 284159:4]
  wire [7:0] d_sizes_clr = _GEN_24[7:0]; // @[chipyard.TestHarness.RocketConfig.fir 284026:4]
  wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56 chipyard.TestHarness.RocketConfig.fir 284160:4]
  wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.RocketConfig.fir 284161:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 284163:4]
  wire  _T_1145 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.RocketConfig.fir 284166:4]
  wire  _T_1146 = ~_T_1145; // @[Monitor.scala 709:16 chipyard.TestHarness.RocketConfig.fir 284167:4]
  wire  _T_1147 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.RocketConfig.fir 284168:4]
  wire  _T_1148 = _T_1146 | _T_1147; // @[Monitor.scala 709:30 chipyard.TestHarness.RocketConfig.fir 284169:4]
  wire  _T_1149 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.RocketConfig.fir 284170:4]
  wire  _T_1150 = _T_1148 | _T_1149; // @[Monitor.scala 709:47 chipyard.TestHarness.RocketConfig.fir 284171:4]
  wire  _T_1152 = _T_1150 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 284173:4]
  wire  _T_1153 = ~_T_1152; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 284174:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.RocketConfig.fir 284180:4]
  wire  _T_1156 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.RocketConfig.fir 284184:4]
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 284190:4]
  reg [8:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 284225:4]
  wire [8:0] d_first_counter1_2 = d_first_counter_2 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 284227:4]
  wire  d_first_2 = d_first_counter_2 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 284228:4]
  wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.RocketConfig.fir 284261:4]
  wire [15:0] _GEN_87 = {{8'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.RocketConfig.fir 284266:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_87 & _a_size_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.RocketConfig.fir 284266:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.RocketConfig.fir 284267:4]
  wire  _T_1174 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.RocketConfig.fir 284345:4]
  wire  _T_1176 = _T_1174 & _T_881; // @[Monitor.scala 779:71 chipyard.TestHarness.RocketConfig.fir 284347:4]
  wire  _T_1178 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.RocketConfig.fir 284353:4]
  wire  _T_1180 = _T_1178 & _T_881; // @[Monitor.scala 783:72 chipyard.TestHarness.RocketConfig.fir 284355:4]
  wire [30:0] _GEN_69 = _T_1180 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.RocketConfig.fir 284356:4 Monitor.scala 786:21 chipyard.TestHarness.RocketConfig.fir 284372:6 chipyard.TestHarness.RocketConfig.fir 284343:4]
  wire  _T_1184 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.RocketConfig.fir 284391:6]
  wire  _T_1188 = _T_1184 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284395:6]
  wire  _T_1189 = ~_T_1188; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284396:6]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.RocketConfig.fir 284249:4 Monitor.scala 747:21 chipyard.TestHarness.RocketConfig.fir 284268:4]
  wire  _T_1194 = _GEN_83 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.RocketConfig.fir 284414:8]
  wire  _T_1196 = _T_1194 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284416:8]
  wire  _T_1197 = ~_T_1196; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284417:8]
  wire [7:0] d_sizes_clr_1 = _GEN_69[7:0]; // @[chipyard.TestHarness.RocketConfig.fir 284342:4]
  wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58 chipyard.TestHarness.RocketConfig.fir 284467:4]
  wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.RocketConfig.fir 284468:4]
  wire  _GEN_93 = io_in_a_valid & _T_15; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282397:10]
  wire  _GEN_109 = io_in_a_valid & _T_171; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282587:10]
  wire  _GEN_127 = io_in_a_valid & _T_331; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282725:10]
  wire  _GEN_141 = io_in_a_valid & _T_426; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282917:10]
  wire  _GEN_151 = io_in_a_valid & _T_517; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283030:10]
  wire  _GEN_161 = io_in_a_valid & _T_610; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283140:10]
  wire  _GEN_171 = io_in_a_valid & _T_696; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283248:10]
  wire  _GEN_181 = io_in_a_valid & _T_782; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283361:10]
  wire  _GEN_193 = io_in_d_valid & _T_881; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283424:10]
  wire  _GEN_203 = io_in_d_valid & _T_901; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283466:10]
  wire  _GEN_213 = io_in_d_valid & _T_929; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283524:10]
  wire  _GEN_223 = io_in_d_valid & _T_958; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283583:10]
  wire  _GEN_229 = io_in_d_valid & _T_975; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283618:10]
  wire  _GEN_235 = io_in_d_valid & _T_993; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283654:10]
  wire  _GEN_241 = _T_1088 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284087:10]
  wire  _GEN_246 = _T_1088 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284109:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 284164:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 284471:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283723:4]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283723:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 283733:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 283734:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 283722:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 283788:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.RocketConfig.fir 283789:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 283788:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.RocketConfig.fir 283790:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 283788:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.RocketConfig.fir 283791:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 283788:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.RocketConfig.fir 283792:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 283788:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.RocketConfig.fir 283793:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283803:4]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283803:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 283813:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 283814:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 283802:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 283877:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.RocketConfig.fir 283878:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 283877:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.RocketConfig.fir 283879:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 283877:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.RocketConfig.fir 283880:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 283877:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.RocketConfig.fir 283881:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 283877:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.RocketConfig.fir 283882:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 283877:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.RocketConfig.fir 283883:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 283885:4]
      inflight <= 1'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 283885:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.RocketConfig.fir 284154:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 283886:4]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 283886:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.RocketConfig.fir 284158:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 283887:4]
      inflight_sizes <= 8'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 283887:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.RocketConfig.fir 284162:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283897:4]
      a_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283897:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 283907:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 283908:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 283722:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 9'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283919:4]
      d_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 283919:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 283929:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 283930:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 283802:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 9'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 284163:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 284163:4]
    end else if (_T_1156) begin // @[Monitor.scala 712:47 chipyard.TestHarness.RocketConfig.fir 284185:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.RocketConfig.fir 284186:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.RocketConfig.fir 284181:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 284190:4]
      inflight_sizes_1 <= 8'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 284190:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.RocketConfig.fir 284469:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 284225:4]
      d_first_counter_2 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 284225:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 284235:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 284236:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 283802:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 9'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_15 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282397:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282398:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282464:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282465:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282471:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282472:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282479:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282480:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282486:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282487:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_161) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282494:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_161) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282495:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282503:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282504:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282511:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282512:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282587:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282588:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282654:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282655:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282661:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282662:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282669:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282670:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282676:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282677:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_161) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282684:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_161) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282685:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_321) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282692:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_321) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282693:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282701:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282702:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282709:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282710:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_331 & _T_340) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282725:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_340) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282726:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_407) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282796:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_407) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282797:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282803:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282804:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282810:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282811:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282818:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282819:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282826:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282827:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282834:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282835:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_426 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282917:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282918:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282924:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282925:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282931:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282932:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282939:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282940:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282947:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 282948:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_517 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283030:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283031:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283037:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283038:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283044:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283045:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283052:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283053:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_609) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283062:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_609) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283063:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_610 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283140:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283141:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283147:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283148:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283154:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283155:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_691) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283162:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_691) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283163:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283170:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283171:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_696 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283248:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283249:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283255:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283256:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283262:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283263:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_777) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283270:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_777) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283271:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283278:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283279:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_782 & _T_858) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283361:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_858) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283362:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283368:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283369:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283375:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283376:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_868) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283383:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_868) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283384:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283391:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283392:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283399:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283400:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283410:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283411:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_881 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283424:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283425:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283432:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283433:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283440:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283441:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283448:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283449:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_900) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283456:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_900) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283457:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_901 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283466:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283467:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283481:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283482:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283489:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283490:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283497:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283498:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283505:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283506:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_929 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283524:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283525:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283539:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283540:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283547:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283548:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283555:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283556:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283564:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283565:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_958 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283583:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283584:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283591:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283592:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283599:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283600:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_975 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283618:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283619:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_229 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283626:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283627:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_229 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283635:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283636:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_993 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283654:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283655:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283662:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283663:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283670:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283671:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283750:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283751:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1031) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283758:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1031) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283759:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283766:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283767:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1039) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283774:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1039) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283775:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283782:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 283783:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283831:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283832:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283839:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283840:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283847:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283848:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283855:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283856:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283863:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283864:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283871:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 283872:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 284016:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 284017:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284076:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284077:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & same_cycle_resp & _T_1109) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284087:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1109) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284088:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1113) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284095:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1113) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284096:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & ~same_cycle_resp & _T_1121) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284109:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_246 & _T_1121) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284110:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_246 & _T_1125) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284117:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_246 & _T_1125) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284118:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284136:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284137:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1144) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 6 (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284148:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1144) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284149:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1153) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 284176:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1153) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 284177:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284398:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284399:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284419:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 284420:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inflight_opcodes = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  inflight_sizes = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_20[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLSerdesser_1_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 284691:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 284692:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 284693:4]
  output        auto_manager_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input         auto_manager_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [2:0]  auto_manager_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [2:0]  auto_manager_in_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [3:0]  auto_manager_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input         auto_manager_in_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [31:0] auto_manager_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [7:0]  auto_manager_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [63:0] auto_manager_in_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input         auto_manager_in_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input         auto_manager_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output        auto_manager_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [2:0]  auto_manager_in_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [1:0]  auto_manager_in_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [3:0]  auto_manager_in_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output        auto_manager_in_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [2:0]  auto_manager_in_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output        auto_manager_in_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [63:0] auto_manager_in_d_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output        auto_manager_in_d_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input         auto_client_out_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output        auto_client_out_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [2:0]  auto_client_out_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [2:0]  auto_client_out_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [2:0]  auto_client_out_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [3:0]  auto_client_out_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [28:0] auto_client_out_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [7:0]  auto_client_out_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output [63:0] auto_client_out_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output        auto_client_out_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output        auto_client_out_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input         auto_client_out_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [2:0]  auto_client_out_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [1:0]  auto_client_out_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [2:0]  auto_client_out_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [3:0]  auto_client_out_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input         auto_client_out_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input         auto_client_out_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input  [63:0] auto_client_out_d_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  input         auto_client_out_d_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 284694:4]
  output        io_ser_in_ready, // @[chipyard.TestHarness.RocketConfig.fir 284695:4]
  input         io_ser_in_valid, // @[chipyard.TestHarness.RocketConfig.fir 284695:4]
  input  [3:0]  io_ser_in_bits, // @[chipyard.TestHarness.RocketConfig.fir 284695:4]
  input         io_ser_out_ready, // @[chipyard.TestHarness.RocketConfig.fir 284695:4]
  output        io_ser_out_valid, // @[chipyard.TestHarness.RocketConfig.fir 284695:4]
  output [3:0]  io_ser_out_bits // @[chipyard.TestHarness.RocketConfig.fir 284695:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire [2:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
  wire  outArb_clock; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_reset; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_in_1_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_in_1_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [2:0] outArb_io_in_1_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [2:0] outArb_io_in_1_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [3:0] outArb_io_in_1_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [3:0] outArb_io_in_1_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [63:0] outArb_io_in_1_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_in_1_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [7:0] outArb_io_in_1_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_in_1_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_in_4_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_in_4_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [2:0] outArb_io_in_4_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [2:0] outArb_io_in_4_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [3:0] outArb_io_in_4_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [3:0] outArb_io_in_4_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [31:0] outArb_io_in_4_bits_address; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [63:0] outArb_io_in_4_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_in_4_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [7:0] outArb_io_in_4_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_in_4_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_out_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_out_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [2:0] outArb_io_out_bits_chanId; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [2:0] outArb_io_out_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [2:0] outArb_io_out_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [3:0] outArb_io_out_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [3:0] outArb_io_out_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [31:0] outArb_io_out_bits_address; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [63:0] outArb_io_out_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_out_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire [7:0] outArb_io_out_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outArb_io_out_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
  wire  outSer_clock; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire  outSer_reset; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire  outSer_io_in_ready; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire  outSer_io_in_valid; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire [2:0] outSer_io_in_bits_chanId; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire [2:0] outSer_io_in_bits_opcode; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire [2:0] outSer_io_in_bits_param; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire [3:0] outSer_io_in_bits_size; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire [3:0] outSer_io_in_bits_source; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire [31:0] outSer_io_in_bits_address; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire [63:0] outSer_io_in_bits_data; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire  outSer_io_in_bits_corrupt; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire [7:0] outSer_io_in_bits_union; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire  outSer_io_in_bits_last; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire  outSer_io_out_ready; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire  outSer_io_out_valid; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire [3:0] outSer_io_out_bits; // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
  wire  inDes_clock; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire  inDes_reset; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire  inDes_io_in_ready; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire  inDes_io_in_valid; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire [3:0] inDes_io_in_bits; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire  inDes_io_out_ready; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire  inDes_io_out_valid; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire [2:0] inDes_io_out_bits_chanId; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire [2:0] inDes_io_out_bits_opcode; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire [2:0] inDes_io_out_bits_param; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire [3:0] inDes_io_out_bits_size; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire [3:0] inDes_io_out_bits_source; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire [31:0] inDes_io_out_bits_address; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire [63:0] inDes_io_out_bits_data; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire  inDes_io_out_bits_corrupt; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire [7:0] inDes_io_out_bits_union; // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
  wire [1:0] _merged_bits_merged_union_T_1 = {auto_client_out_d_bits_sink,auto_client_out_d_bits_denied}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 284794:4]
  wire  merged_1_ready = outArb_io_in_1_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.RocketConfig.fir 284783:4 Serdes.scala 625:18 chipyard.TestHarness.RocketConfig.fir 284979:4]
  wire  _merged_bits_last_T_1 = merged_1_ready & auto_client_out_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 284807:4]
  wire [12:0] _merged_bits_last_beats1_decode_T_1 = 13'h3f << auto_client_out_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 284809:4]
  wire [5:0] _merged_bits_last_beats1_decode_T_3 = ~_merged_bits_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 284811:4]
  wire [2:0] merged_bits_last_beats1_decode = _merged_bits_last_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.RocketConfig.fir 284812:4]
  wire  merged_bits_last_beats1_opdata = auto_client_out_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.RocketConfig.fir 284813:4]
  wire [2:0] merged_bits_last_beats1 = merged_bits_last_beats1_opdata ? merged_bits_last_beats1_decode : 3'h0; // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 284814:4]
  reg [2:0] merged_bits_last_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 284815:4]
  wire [2:0] merged_bits_last_counter1_1 = merged_bits_last_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 284817:4]
  wire  merged_bits_last_first_1 = merged_bits_last_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 284818:4]
  wire  _merged_bits_last_last_T_2 = merged_bits_last_counter_1 == 3'h1; // @[Edges.scala 231:25 chipyard.TestHarness.RocketConfig.fir 284819:4]
  wire  _merged_bits_last_last_T_3 = merged_bits_last_beats1 == 3'h0; // @[Edges.scala 231:47 chipyard.TestHarness.RocketConfig.fir 284820:4]
  wire  merged_4_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.RocketConfig.fir 284926:4 Serdes.scala 625:18 chipyard.TestHarness.RocketConfig.fir 284988:4]
  wire  _merged_bits_last_T_4 = merged_4_ready & auto_manager_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 284949:4]
  wire [20:0] _merged_bits_last_beats1_decode_T_13 = 21'h3f << auto_manager_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 284951:4]
  wire [5:0] _merged_bits_last_beats1_decode_T_15 = ~_merged_bits_last_beats1_decode_T_13[5:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 284953:4]
  wire [2:0] merged_bits_last_beats1_decode_3 = _merged_bits_last_beats1_decode_T_15[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.RocketConfig.fir 284954:4]
  wire  merged_bits_last_beats1_opdata_3 = ~auto_manager_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.RocketConfig.fir 284956:4]
  wire [2:0] merged_bits_last_beats1_3 = merged_bits_last_beats1_opdata_3 ? merged_bits_last_beats1_decode_3 : 3'h0; // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 284957:4]
  reg [2:0] merged_bits_last_counter_4; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 284958:4]
  wire [2:0] merged_bits_last_counter1_4 = merged_bits_last_counter_4 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 284960:4]
  wire  merged_bits_last_first_4 = merged_bits_last_counter_4 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 284961:4]
  wire  _merged_bits_last_last_T_8 = merged_bits_last_counter_4 == 3'h1; // @[Edges.scala 231:25 chipyard.TestHarness.RocketConfig.fir 284962:4]
  wire  _merged_bits_last_last_T_9 = merged_bits_last_beats1_3 == 3'h0; // @[Edges.scala 231:47 chipyard.TestHarness.RocketConfig.fir 284963:4]
  wire  _bundleOut_0_a_valid_T = inDes_io_out_bits_chanId == 3'h0; // @[Serdes.scala 236:37 chipyard.TestHarness.RocketConfig.fir 285001:4]
  wire  _bundleIn_0_d_valid_T = inDes_io_out_bits_chanId == 3'h3; // @[Serdes.scala 239:37 chipyard.TestHarness.RocketConfig.fir 285067:4]
  wire [7:0] _bundleIn_0_d_bits_d_sink_T = {{1'd0}, inDes_io_out_bits_union[7:1]}; // @[Serdes.scala 468:31 chipyard.TestHarness.RocketConfig.fir 285077:4]
  wire  _inDes_io_out_ready_T = 3'h0 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.RocketConfig.fir 285106:4]
  wire  _inDes_io_out_ready_T_1 = _inDes_io_out_ready_T & auto_client_out_a_ready; // @[Mux.scala 80:57 chipyard.TestHarness.RocketConfig.fir 285107:4]
  wire  _inDes_io_out_ready_T_2 = 3'h1 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.RocketConfig.fir 285108:4]
  wire  _inDes_io_out_ready_T_3 = _inDes_io_out_ready_T_2 ? 1'h0 : _inDes_io_out_ready_T_1; // @[Mux.scala 80:57 chipyard.TestHarness.RocketConfig.fir 285109:4]
  wire  _inDes_io_out_ready_T_4 = 3'h2 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.RocketConfig.fir 285110:4]
  wire  _inDes_io_out_ready_T_5 = _inDes_io_out_ready_T_4 ? 1'h0 : _inDes_io_out_ready_T_3; // @[Mux.scala 80:57 chipyard.TestHarness.RocketConfig.fir 285111:4]
  wire  _inDes_io_out_ready_T_6 = 3'h3 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.RocketConfig.fir 285112:4]
  wire  _inDes_io_out_ready_T_7 = _inDes_io_out_ready_T_6 ? auto_manager_in_d_ready : _inDes_io_out_ready_T_5; // @[Mux.scala 80:57 chipyard.TestHarness.RocketConfig.fir 285113:4]
  wire  _inDes_io_out_ready_T_8 = 3'h4 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.RocketConfig.fir 285114:4]
  TLMonitor_53_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 284705:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  HellaPeekingArbiter_inTestHarness outArb ( // @[Serdes.scala 622:24 chipyard.TestHarness.RocketConfig.fir 284736:4]
    .clock(outArb_clock),
    .reset(outArb_reset),
    .io_in_1_ready(outArb_io_in_1_ready),
    .io_in_1_valid(outArb_io_in_1_valid),
    .io_in_1_bits_opcode(outArb_io_in_1_bits_opcode),
    .io_in_1_bits_param(outArb_io_in_1_bits_param),
    .io_in_1_bits_size(outArb_io_in_1_bits_size),
    .io_in_1_bits_source(outArb_io_in_1_bits_source),
    .io_in_1_bits_data(outArb_io_in_1_bits_data),
    .io_in_1_bits_corrupt(outArb_io_in_1_bits_corrupt),
    .io_in_1_bits_union(outArb_io_in_1_bits_union),
    .io_in_1_bits_last(outArb_io_in_1_bits_last),
    .io_in_4_ready(outArb_io_in_4_ready),
    .io_in_4_valid(outArb_io_in_4_valid),
    .io_in_4_bits_opcode(outArb_io_in_4_bits_opcode),
    .io_in_4_bits_param(outArb_io_in_4_bits_param),
    .io_in_4_bits_size(outArb_io_in_4_bits_size),
    .io_in_4_bits_source(outArb_io_in_4_bits_source),
    .io_in_4_bits_address(outArb_io_in_4_bits_address),
    .io_in_4_bits_data(outArb_io_in_4_bits_data),
    .io_in_4_bits_corrupt(outArb_io_in_4_bits_corrupt),
    .io_in_4_bits_union(outArb_io_in_4_bits_union),
    .io_in_4_bits_last(outArb_io_in_4_bits_last),
    .io_out_ready(outArb_io_out_ready),
    .io_out_valid(outArb_io_out_valid),
    .io_out_bits_chanId(outArb_io_out_bits_chanId),
    .io_out_bits_opcode(outArb_io_out_bits_opcode),
    .io_out_bits_param(outArb_io_out_bits_param),
    .io_out_bits_size(outArb_io_out_bits_size),
    .io_out_bits_source(outArb_io_out_bits_source),
    .io_out_bits_address(outArb_io_out_bits_address),
    .io_out_bits_data(outArb_io_out_bits_data),
    .io_out_bits_corrupt(outArb_io_out_bits_corrupt),
    .io_out_bits_union(outArb_io_out_bits_union),
    .io_out_bits_last(outArb_io_out_bits_last)
  );
  GenericSerializer_inTestHarness outSer ( // @[Serdes.scala 624:24 chipyard.TestHarness.RocketConfig.fir 284739:4]
    .clock(outSer_clock),
    .reset(outSer_reset),
    .io_in_ready(outSer_io_in_ready),
    .io_in_valid(outSer_io_in_valid),
    .io_in_bits_chanId(outSer_io_in_bits_chanId),
    .io_in_bits_opcode(outSer_io_in_bits_opcode),
    .io_in_bits_param(outSer_io_in_bits_param),
    .io_in_bits_size(outSer_io_in_bits_size),
    .io_in_bits_source(outSer_io_in_bits_source),
    .io_in_bits_address(outSer_io_in_bits_address),
    .io_in_bits_data(outSer_io_in_bits_data),
    .io_in_bits_corrupt(outSer_io_in_bits_corrupt),
    .io_in_bits_union(outSer_io_in_bits_union),
    .io_in_bits_last(outSer_io_in_bits_last),
    .io_out_ready(outSer_io_out_ready),
    .io_out_valid(outSer_io_out_valid),
    .io_out_bits(outSer_io_out_bits)
  );
  GenericDeserializer_inTestHarness inDes ( // @[Serdes.scala 629:23 chipyard.TestHarness.RocketConfig.fir 284995:4]
    .clock(inDes_clock),
    .reset(inDes_reset),
    .io_in_ready(inDes_io_in_ready),
    .io_in_valid(inDes_io_in_valid),
    .io_in_bits(inDes_io_in_bits),
    .io_out_ready(inDes_io_out_ready),
    .io_out_valid(inDes_io_out_valid),
    .io_out_bits_chanId(inDes_io_out_bits_chanId),
    .io_out_bits_opcode(inDes_io_out_bits_opcode),
    .io_out_bits_param(inDes_io_out_bits_param),
    .io_out_bits_size(inDes_io_out_bits_size),
    .io_out_bits_source(inDes_io_out_bits_source),
    .io_out_bits_address(inDes_io_out_bits_address),
    .io_out_bits_data(inDes_io_out_bits_data),
    .io_out_bits_corrupt(inDes_io_out_bits_corrupt),
    .io_out_bits_union(inDes_io_out_bits_union)
  );
  assign auto_manager_in_a_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.RocketConfig.fir 284926:4 Serdes.scala 625:18 chipyard.TestHarness.RocketConfig.fir 284988:4]
  assign auto_manager_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 637:46 chipyard.TestHarness.RocketConfig.fir 285068:4]
  assign auto_manager_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 461:15 chipyard.TestHarness.RocketConfig.fir 285071:4]
  assign auto_manager_in_d_bits_param = inDes_io_out_bits_param[1:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 462:15 chipyard.TestHarness.RocketConfig.fir 285072:4]
  assign auto_manager_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 463:15 chipyard.TestHarness.RocketConfig.fir 285073:4]
  assign auto_manager_in_d_bits_source = inDes_io_out_bits_source[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 464:15 chipyard.TestHarness.RocketConfig.fir 285074:4]
  assign auto_manager_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[2:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 468:17 chipyard.TestHarness.RocketConfig.fir 285078:4]
  assign auto_manager_in_d_bits_denied = inDes_io_out_bits_union[0]; // @[Serdes.scala 469:30 chipyard.TestHarness.RocketConfig.fir 285079:4]
  assign auto_manager_in_d_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 465:15 chipyard.TestHarness.RocketConfig.fir 285075:4]
  assign auto_manager_in_d_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 467:17 chipyard.TestHarness.RocketConfig.fir 285076:4]
  assign auto_client_out_a_valid = inDes_io_out_valid & _bundleOut_0_a_valid_T; // @[Serdes.scala 631:45 chipyard.TestHarness.RocketConfig.fir 285002:4]
  assign auto_client_out_a_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 374:17 chipyard.TestHarness.RocketConfig.fir 285004:4 Serdes.scala 375:15 chipyard.TestHarness.RocketConfig.fir 285005:4]
  assign auto_client_out_a_bits_param = inDes_io_out_bits_param; // @[Serdes.scala 374:17 chipyard.TestHarness.RocketConfig.fir 285004:4 Serdes.scala 376:15 chipyard.TestHarness.RocketConfig.fir 285006:4]
  assign auto_client_out_a_bits_size = inDes_io_out_bits_size[2:0]; // @[Serdes.scala 374:17 chipyard.TestHarness.RocketConfig.fir 285004:4 Serdes.scala 377:15 chipyard.TestHarness.RocketConfig.fir 285007:4]
  assign auto_client_out_a_bits_source = inDes_io_out_bits_source; // @[Serdes.scala 374:17 chipyard.TestHarness.RocketConfig.fir 285004:4 Serdes.scala 378:15 chipyard.TestHarness.RocketConfig.fir 285008:4]
  assign auto_client_out_a_bits_address = inDes_io_out_bits_address[28:0]; // @[Serdes.scala 374:17 chipyard.TestHarness.RocketConfig.fir 285004:4 Serdes.scala 379:15 chipyard.TestHarness.RocketConfig.fir 285009:4]
  assign auto_client_out_a_bits_mask = inDes_io_out_bits_union; // @[Serdes.scala 374:17 chipyard.TestHarness.RocketConfig.fir 285004:4 Serdes.scala 385:15 chipyard.TestHarness.RocketConfig.fir 285012:4]
  assign auto_client_out_a_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 374:17 chipyard.TestHarness.RocketConfig.fir 285004:4 Serdes.scala 380:15 chipyard.TestHarness.RocketConfig.fir 285010:4]
  assign auto_client_out_a_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 374:17 chipyard.TestHarness.RocketConfig.fir 285004:4 Serdes.scala 382:17 chipyard.TestHarness.RocketConfig.fir 285011:4]
  assign auto_client_out_d_ready = outArb_io_in_1_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.RocketConfig.fir 284783:4 Serdes.scala 625:18 chipyard.TestHarness.RocketConfig.fir 284979:4]
  assign io_ser_in_ready = inDes_io_in_ready; // @[Serdes.scala 630:17 chipyard.TestHarness.RocketConfig.fir 285000:4]
  assign io_ser_out_valid = outSer_io_out_valid; // @[Serdes.scala 627:16 chipyard.TestHarness.RocketConfig.fir 284993:4]
  assign io_ser_out_bits = outSer_io_out_bits; // @[Serdes.scala 627:16 chipyard.TestHarness.RocketConfig.fir 284992:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 284706:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 284707:4]
  assign monitor_io_in_a_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.RocketConfig.fir 284926:4 Serdes.scala 625:18 chipyard.TestHarness.RocketConfig.fir 284988:4]
  assign monitor_io_in_a_valid = auto_manager_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign monitor_io_in_a_bits_opcode = auto_manager_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign monitor_io_in_a_bits_param = auto_manager_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign monitor_io_in_a_bits_size = auto_manager_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign monitor_io_in_a_bits_source = auto_manager_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign monitor_io_in_a_bits_address = auto_manager_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign monitor_io_in_a_bits_mask = auto_manager_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign monitor_io_in_a_bits_corrupt = auto_manager_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign monitor_io_in_d_ready = auto_manager_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign monitor_io_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 637:46 chipyard.TestHarness.RocketConfig.fir 285068:4]
  assign monitor_io_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 461:15 chipyard.TestHarness.RocketConfig.fir 285071:4]
  assign monitor_io_in_d_bits_param = inDes_io_out_bits_param[1:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 462:15 chipyard.TestHarness.RocketConfig.fir 285072:4]
  assign monitor_io_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 463:15 chipyard.TestHarness.RocketConfig.fir 285073:4]
  assign monitor_io_in_d_bits_source = inDes_io_out_bits_source[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 464:15 chipyard.TestHarness.RocketConfig.fir 285074:4]
  assign monitor_io_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[2:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 468:17 chipyard.TestHarness.RocketConfig.fir 285078:4]
  assign monitor_io_in_d_bits_denied = inDes_io_out_bits_union[0]; // @[Serdes.scala 469:30 chipyard.TestHarness.RocketConfig.fir 285079:4]
  assign monitor_io_in_d_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 460:17 chipyard.TestHarness.RocketConfig.fir 285070:4 Serdes.scala 467:17 chipyard.TestHarness.RocketConfig.fir 285076:4]
  assign outArb_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 284737:4]
  assign outArb_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 284738:4]
  assign outArb_io_in_1_valid = auto_client_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 284701:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 284728:4]
  assign outArb_io_in_1_bits_opcode = auto_client_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 284701:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 284728:4]
  assign outArb_io_in_1_bits_param = {{1'd0}, auto_client_out_d_bits_param}; // @[Serdes.scala 312:22 chipyard.TestHarness.RocketConfig.fir 284785:4 Serdes.scala 315:20 chipyard.TestHarness.RocketConfig.fir 284788:4]
  assign outArb_io_in_1_bits_size = {{1'd0}, auto_client_out_d_bits_size}; // @[Serdes.scala 312:22 chipyard.TestHarness.RocketConfig.fir 284785:4 Serdes.scala 316:20 chipyard.TestHarness.RocketConfig.fir 284789:4]
  assign outArb_io_in_1_bits_source = auto_client_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 284701:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 284728:4]
  assign outArb_io_in_1_bits_data = auto_client_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 284701:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 284728:4]
  assign outArb_io_in_1_bits_corrupt = auto_client_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 284701:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 284728:4]
  assign outArb_io_in_1_bits_union = {{6'd0}, _merged_bits_merged_union_T_1}; // @[Serdes.scala 312:22 chipyard.TestHarness.RocketConfig.fir 284785:4 Serdes.scala 322:22 chipyard.TestHarness.RocketConfig.fir 284795:4]
  assign outArb_io_in_1_bits_last = _merged_bits_last_last_T_2 | _merged_bits_last_last_T_3; // @[Edges.scala 231:37 chipyard.TestHarness.RocketConfig.fir 284821:4]
  assign outArb_io_in_4_valid = auto_manager_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign outArb_io_in_4_bits_opcode = auto_manager_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign outArb_io_in_4_bits_param = auto_manager_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign outArb_io_in_4_bits_size = auto_manager_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign outArb_io_in_4_bits_source = {{3'd0}, auto_manager_in_a_bits_source}; // @[Serdes.scala 255:22 chipyard.TestHarness.RocketConfig.fir 284928:4 Serdes.scala 260:20 chipyard.TestHarness.RocketConfig.fir 284933:4]
  assign outArb_io_in_4_bits_address = auto_manager_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign outArb_io_in_4_bits_data = auto_manager_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign outArb_io_in_4_bits_corrupt = auto_manager_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign outArb_io_in_4_bits_union = auto_manager_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 284703:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 284729:4]
  assign outArb_io_in_4_bits_last = _merged_bits_last_last_T_8 | _merged_bits_last_last_T_9; // @[Edges.scala 231:37 chipyard.TestHarness.RocketConfig.fir 284964:4]
  assign outArb_io_out_ready = outSer_io_in_ready; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284991:4]
  assign outSer_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 284740:4]
  assign outSer_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 284741:4]
  assign outSer_io_in_valid = outArb_io_out_valid; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284990:4]
  assign outSer_io_in_bits_chanId = outArb_io_out_bits_chanId; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284989:4]
  assign outSer_io_in_bits_opcode = outArb_io_out_bits_opcode; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284989:4]
  assign outSer_io_in_bits_param = outArb_io_out_bits_param; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284989:4]
  assign outSer_io_in_bits_size = outArb_io_out_bits_size; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284989:4]
  assign outSer_io_in_bits_source = outArb_io_out_bits_source; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284989:4]
  assign outSer_io_in_bits_address = outArb_io_out_bits_address; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284989:4]
  assign outSer_io_in_bits_data = outArb_io_out_bits_data; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284989:4]
  assign outSer_io_in_bits_corrupt = outArb_io_out_bits_corrupt; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284989:4]
  assign outSer_io_in_bits_union = outArb_io_out_bits_union; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284989:4]
  assign outSer_io_in_bits_last = outArb_io_out_bits_last; // @[Serdes.scala 626:18 chipyard.TestHarness.RocketConfig.fir 284989:4]
  assign outSer_io_out_ready = io_ser_out_ready; // @[Serdes.scala 627:16 chipyard.TestHarness.RocketConfig.fir 284994:4]
  assign inDes_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 284996:4]
  assign inDes_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 284997:4]
  assign inDes_io_in_valid = io_ser_in_valid; // @[Serdes.scala 630:17 chipyard.TestHarness.RocketConfig.fir 284999:4]
  assign inDes_io_in_bits = io_ser_in_bits; // @[Serdes.scala 630:17 chipyard.TestHarness.RocketConfig.fir 284998:4]
  assign inDes_io_out_ready = _inDes_io_out_ready_T_8 ? 1'h0 : _inDes_io_out_ready_T_7; // @[Mux.scala 80:57 chipyard.TestHarness.RocketConfig.fir 285115:4]
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 284815:4]
      merged_bits_last_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 284815:4]
    end else if (_merged_bits_last_T_1) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 284825:4]
      if (merged_bits_last_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 284826:6]
        if (merged_bits_last_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 284814:4]
          merged_bits_last_counter_1 <= merged_bits_last_beats1_decode;
        end else begin
          merged_bits_last_counter_1 <= 3'h0;
        end
      end else begin
        merged_bits_last_counter_1 <= merged_bits_last_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 284958:4]
      merged_bits_last_counter_4 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 284958:4]
    end else if (_merged_bits_last_T_4) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 284968:4]
      if (merged_bits_last_first_4) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 284969:6]
        if (merged_bits_last_beats1_opdata_3) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 284957:4]
          merged_bits_last_counter_4 <= merged_bits_last_beats1_decode_3;
        end else begin
          merged_bits_last_counter_4 <= 3'h0;
        end
      end else begin
        merged_bits_last_counter_4 <= merged_bits_last_counter1_4;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  merged_bits_last_counter_1 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  merged_bits_last_counter_4 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_54_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 285134:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 285135:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 285136:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input  [1:0]  io_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input  [7:0]  io_in_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input  [1:0]  io_in_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
  input  [7:0]  io_in_d_bits_source // @[chipyard.TestHarness.RocketConfig.fir 285137:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [159:0] _RAND_10;
  reg [639:0] _RAND_11;
  reg [639:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [159:0] _RAND_16;
  reg [639:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 286628:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 286935:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.RocketConfig.fir 285154:6]
  wire [5:0] _is_aligned_mask_T_1 = 6'h7 << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 285160:6]
  wire [2:0] is_aligned_mask = ~_is_aligned_mask_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 285162:6]
  wire [28:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.RocketConfig.fir 285163:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.RocketConfig.fir 285163:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.RocketConfig.fir 285164:6]
  wire [2:0] _mask_sizeOH_T = {{1'd0}, io_in_a_bits_size}; // @[Misc.scala 201:34 chipyard.TestHarness.RocketConfig.fir 285165:6]
  wire [1:0] mask_sizeOH_shiftAmount = _mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.RocketConfig.fir 285166:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.RocketConfig.fir 285167:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.RocketConfig.fir 285169:6]
  wire  _mask_T = io_in_a_bits_size >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.RocketConfig.fir 285170:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 285171:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 285172:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 285173:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285175:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285176:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285178:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285179:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 285180:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 285181:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 285182:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285183:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285184:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285185:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285186:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285187:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285188:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285189:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285190:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285191:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285192:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285193:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285194:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 285195:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 285196:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 285197:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285198:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285199:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285200:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285201:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285202:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285203:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285204:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285205:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285206:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285207:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285208:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285209:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285210:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285211:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285212:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285213:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285214:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285215:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285216:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285217:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285218:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 285219:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 285220:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 285221:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 285228:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.RocketConfig.fir 285251:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 285267:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 285268:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 285270:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 285271:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285277:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285302:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285303:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285310:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285311:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285317:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285318:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.RocketConfig.fir 285323:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285325:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285326:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.RocketConfig.fir 285331:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.RocketConfig.fir 285332:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285334:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285335:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.RocketConfig.fir 285340:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285342:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285343:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.RocketConfig.fir 285349:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.RocketConfig.fir 285429:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285431:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285432:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.RocketConfig.fir 285455:6]
  wire  _T_175 = _T_37 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285489:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285490:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.RocketConfig.fir 285509:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285511:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285512:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.RocketConfig.fir 285517:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285519:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285520:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.RocketConfig.fir 285534:6]
  wire  _T_218 = _source_ok_T_4 & _T_37; // @[Monitor.scala 115:71 chipyard.TestHarness.RocketConfig.fir 285560:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285562:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285563:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.RocketConfig.fir 285599:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.RocketConfig.fir 285655:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.RocketConfig.fir 285656:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.RocketConfig.fir 285657:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285659:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285660:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.RocketConfig.fir 285666:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.RocketConfig.fir 285711:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285713:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285714:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.RocketConfig.fir 285728:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.RocketConfig.fir 285773:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285775:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285776:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.RocketConfig.fir 285790:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.RocketConfig.fir 285835:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285837:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285838:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.RocketConfig.fir 285862:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285864:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285865:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.RocketConfig.fir 285876:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.RocketConfig.fir 285882:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285885:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285886:8]
  wire  _T_405 = io_in_d_bits_size >= 2'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.RocketConfig.fir 285891:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285893:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285894:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.RocketConfig.fir 285924:6]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.RocketConfig.fir 285982:6]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.RocketConfig.fir 286041:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.RocketConfig.fir 286076:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.RocketConfig.fir 286112:6]
  wire  a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 286178:4]
  reg  a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286187:4]
  wire  a_first_counter1 = a_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 286189:4]
  wire  a_first = ~a_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 286190:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.RocketConfig.fir 286201:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.RocketConfig.fir 286202:4]
  reg [1:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.RocketConfig.fir 286203:4]
  reg [7:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.RocketConfig.fir 286204:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.RocketConfig.fir 286205:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.RocketConfig.fir 286206:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.RocketConfig.fir 286207:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.RocketConfig.fir 286209:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286211:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286212:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.RocketConfig.fir 286217:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286219:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286220:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.RocketConfig.fir 286225:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286227:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286228:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.RocketConfig.fir 286233:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286235:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286236:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.RocketConfig.fir 286241:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286243:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286244:6]
  wire  _T_565 = a_first_done & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.RocketConfig.fir 286251:4]
  wire  d_first_done = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 286259:4]
  reg  d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286267:4]
  wire  d_first_counter1 = d_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 286269:4]
  wire  d_first = ~d_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 286270:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.RocketConfig.fir 286281:4]
  reg [1:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.RocketConfig.fir 286283:4]
  reg [7:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.RocketConfig.fir 286284:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.RocketConfig.fir 286287:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.RocketConfig.fir 286288:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.RocketConfig.fir 286290:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286292:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286293:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.RocketConfig.fir 286306:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286308:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286309:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.RocketConfig.fir 286314:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286316:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286317:6]
  wire  _T_593 = d_first_done & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.RocketConfig.fir 286340:4]
  reg [159:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 286349:4]
  reg [639:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 286350:4]
  reg [639:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 286351:4]
  reg  a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286361:4]
  wire  a_first_counter1_1 = a_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 286363:4]
  wire  a_first_1 = ~a_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 286364:4]
  reg  d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286383:4]
  wire  d_first_counter1_1 = d_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 286385:4]
  wire  d_first_1 = ~d_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 286386:4]
  wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.RocketConfig.fir 286407:4]
  wire [10:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.RocketConfig.fir 286407:4]
  wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.RocketConfig.fir 286408:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.RocketConfig.fir 286412:4]
  wire [639:0] _GEN_73 = {{624'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.RocketConfig.fir 286413:4]
  wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.RocketConfig.fir 286413:4]
  wire [639:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[639:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.RocketConfig.fir 286414:4]
  wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.RocketConfig.fir 286419:4]
  wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.RocketConfig.fir 286424:4]
  wire [639:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[639:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.RocketConfig.fir 286425:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.RocketConfig.fir 286449:4]
  wire [255:0] _a_set_wo_ready_T = 256'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.RocketConfig.fir 286452:6]
  wire [255:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.RocketConfig.fir 286451:4 Monitor.scala 649:22 chipyard.TestHarness.RocketConfig.fir 286453:6 chipyard.TestHarness.RocketConfig.fir 286400:4]
  wire  _T_597 = a_first_done & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.RocketConfig.fir 286456:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.RocketConfig.fir 286461:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.RocketConfig.fir 286462:6]
  wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.RocketConfig.fir 286464:6]
  wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.RocketConfig.fir 286465:6]
  wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.RocketConfig.fir 286467:6]
  wire [10:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.RocketConfig.fir 286467:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 286458:4 Monitor.scala 654:28 chipyard.TestHarness.RocketConfig.fir 286463:6 chipyard.TestHarness.RocketConfig.fir 286446:4]
  wire [2050:0] _GEN_79 = {{2047'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.RocketConfig.fir 286468:6]
  wire [2050:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.RocketConfig.fir 286468:6]
  wire [2:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 3'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 286458:4 Monitor.scala 655:28 chipyard.TestHarness.RocketConfig.fir 286466:6 chipyard.TestHarness.RocketConfig.fir 286448:4]
  wire [2049:0] _GEN_81 = {{2047'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.RocketConfig.fir 286471:6]
  wire [2049:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.RocketConfig.fir 286471:6]
  wire [159:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.RocketConfig.fir 286473:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.RocketConfig.fir 286475:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286477:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286478:6]
  wire [255:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 286458:4 Monitor.scala 653:28 chipyard.TestHarness.RocketConfig.fir 286460:6 chipyard.TestHarness.RocketConfig.fir 286398:4]
  wire [2050:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 2051'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 286458:4 Monitor.scala 656:28 chipyard.TestHarness.RocketConfig.fir 286469:6 chipyard.TestHarness.RocketConfig.fir 286402:4]
  wire [2049:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 2050'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 286458:4 Monitor.scala 657:28 chipyard.TestHarness.RocketConfig.fir 286472:6 chipyard.TestHarness.RocketConfig.fir 286404:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.RocketConfig.fir 286493:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.RocketConfig.fir 286495:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.RocketConfig.fir 286496:4]
  wire [255:0] _d_clr_wo_ready_T = 256'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.RocketConfig.fir 286498:6]
  wire [255:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.RocketConfig.fir 286497:4 Monitor.scala 672:22 chipyard.TestHarness.RocketConfig.fir 286499:6 chipyard.TestHarness.RocketConfig.fir 286487:4]
  wire  _T_610 = d_first_done & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.RocketConfig.fir 286502:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.RocketConfig.fir 286505:4]
  wire [2062:0] _GEN_83 = {{2047'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.RocketConfig.fir 286514:6]
  wire [2062:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.RocketConfig.fir 286514:6]
  wire [255:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 286506:4 Monitor.scala 676:21 chipyard.TestHarness.RocketConfig.fir 286508:6 chipyard.TestHarness.RocketConfig.fir 286485:4]
  wire [2062:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 286506:4 Monitor.scala 677:21 chipyard.TestHarness.RocketConfig.fir 286515:6 chipyard.TestHarness.RocketConfig.fir 286489:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.RocketConfig.fir 286531:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.RocketConfig.fir 286532:6]
  wire [159:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.RocketConfig.fir 286533:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.RocketConfig.fir 286535:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286537:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286538:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 286544:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 286545:8 Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 286545:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 286545:8 Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 286545:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 286545:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.RocketConfig.fir 286546:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286548:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286549:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.RocketConfig.fir 286554:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286556:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286557:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 286405:4 Monitor.scala 634:21 chipyard.TestHarness.RocketConfig.fir 286415:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 286565:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 286567:8 Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 286567:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 286567:8 Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 286567:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 286567:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.RocketConfig.fir 286568:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286570:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286571:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 286416:4 Monitor.scala 638:19 chipyard.TestHarness.RocketConfig.fir 286426:4]
  wire [3:0] _GEN_86 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.RocketConfig.fir 286576:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.RocketConfig.fir 286576:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286578:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286579:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.RocketConfig.fir 286587:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.RocketConfig.fir 286588:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.RocketConfig.fir 286590:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.RocketConfig.fir 286592:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.RocketConfig.fir 286594:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.RocketConfig.fir 286595:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286597:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286598:6]
  wire [159:0] a_set_wo_ready = _GEN_15[159:0]; // @[chipyard.TestHarness.RocketConfig.fir 286399:4]
  wire [159:0] d_clr_wo_ready = _GEN_21[159:0]; // @[chipyard.TestHarness.RocketConfig.fir 286486:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.RocketConfig.fir 286604:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.RocketConfig.fir 286605:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.RocketConfig.fir 286606:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.RocketConfig.fir 286607:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286609:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286610:4]
  wire [159:0] a_set = _GEN_16[159:0]; // @[chipyard.TestHarness.RocketConfig.fir 286397:4]
  wire [159:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.RocketConfig.fir 286615:4]
  wire [159:0] d_clr = _GEN_22[159:0]; // @[chipyard.TestHarness.RocketConfig.fir 286484:4]
  wire [159:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.RocketConfig.fir 286616:4]
  wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.RocketConfig.fir 286617:4]
  wire [639:0] a_opcodes_set = _GEN_19[639:0]; // @[chipyard.TestHarness.RocketConfig.fir 286401:4]
  wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.RocketConfig.fir 286619:4]
  wire [639:0] d_opcodes_clr = _GEN_23[639:0]; // @[chipyard.TestHarness.RocketConfig.fir 286488:4]
  wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.RocketConfig.fir 286620:4]
  wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.RocketConfig.fir 286621:4]
  wire [639:0] a_sizes_set = _GEN_20[639:0]; // @[chipyard.TestHarness.RocketConfig.fir 286403:4]
  wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.RocketConfig.fir 286623:4]
  wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.RocketConfig.fir 286625:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 286627:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.RocketConfig.fir 286630:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.RocketConfig.fir 286631:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.RocketConfig.fir 286632:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.RocketConfig.fir 286633:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.RocketConfig.fir 286634:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.RocketConfig.fir 286635:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286637:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286638:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.RocketConfig.fir 286644:4]
  wire  _T_676 = a_first_done | d_first_done; // @[Monitor.scala 712:27 chipyard.TestHarness.RocketConfig.fir 286648:4]
  reg [159:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.RocketConfig.fir 286652:4]
  reg [639:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 286654:4]
  reg  d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286689:4]
  wire  d_first_counter1_2 = d_first_counter_2 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 286691:4]
  wire  d_first_2 = ~d_first_counter_2; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 286692:4]
  wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.RocketConfig.fir 286725:4]
  wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.RocketConfig.fir 286730:4]
  wire [639:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[639:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.RocketConfig.fir 286731:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.RocketConfig.fir 286809:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.RocketConfig.fir 286811:4]
  wire  _T_698 = d_first_done & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.RocketConfig.fir 286817:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.RocketConfig.fir 286819:4]
  wire [255:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.RocketConfig.fir 286820:4 Monitor.scala 784:21 chipyard.TestHarness.RocketConfig.fir 286822:6 chipyard.TestHarness.RocketConfig.fir 286801:4]
  wire [2062:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.RocketConfig.fir 286820:4 Monitor.scala 785:21 chipyard.TestHarness.RocketConfig.fir 286829:6 chipyard.TestHarness.RocketConfig.fir 286805:4]
  wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.RocketConfig.fir 286855:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286859:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286860:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 286713:4 Monitor.scala 747:21 chipyard.TestHarness.RocketConfig.fir 286732:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.RocketConfig.fir 286878:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286880:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286881:8]
  wire [159:0] d_clr_1 = _GEN_67[159:0]; // @[chipyard.TestHarness.RocketConfig.fir 286800:4]
  wire [159:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.RocketConfig.fir 286923:4]
  wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.RocketConfig.fir 286924:4]
  wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0]; // @[chipyard.TestHarness.RocketConfig.fir 286804:4]
  wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.RocketConfig.fir 286927:4]
  wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.RocketConfig.fir 286932:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.RocketConfig.fir 286934:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.RocketConfig.fir 286937:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.RocketConfig.fir 286938:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.RocketConfig.fir 286939:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.RocketConfig.fir 286940:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.RocketConfig.fir 286941:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.RocketConfig.fir 286942:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286944:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286945:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.RocketConfig.fir 286951:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285279:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285377:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285474:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285565:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285630:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285694:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285756:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285818:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285888:10]
  wire  _GEN_202 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285930:10]
  wire  _GEN_208 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285988:10]
  wire  _GEN_214 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286047:10]
  wire  _GEN_216 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286082:10]
  wire  _GEN_218 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286118:10]
  wire  _GEN_220 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286551:10]
  wire  _GEN_225 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286573:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 286628:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 286935:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286187:4]
      a_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286187:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 286197:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 286198:6]
        a_first_counter <= 1'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 286252:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.RocketConfig.fir 286253:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 286252:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.RocketConfig.fir 286254:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 286252:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.RocketConfig.fir 286255:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 286252:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.RocketConfig.fir 286256:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 286252:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.RocketConfig.fir 286257:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286267:4]
      d_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286267:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 286277:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 286278:6]
        d_first_counter <= 1'h0;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 286341:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.RocketConfig.fir 286342:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 286341:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.RocketConfig.fir 286344:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 286341:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.RocketConfig.fir 286345:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 286349:4]
      inflight <= 160'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 286349:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.RocketConfig.fir 286618:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 286350:4]
      inflight_opcodes <= 640'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 286350:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.RocketConfig.fir 286622:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 286351:4]
      inflight_sizes <= 640'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 286351:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.RocketConfig.fir 286626:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286361:4]
      a_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286361:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 286371:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 286372:6]
        a_first_counter_1 <= 1'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286383:4]
      d_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286383:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 286393:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 286394:6]
        d_first_counter_1 <= 1'h0;
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 286627:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 286627:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.RocketConfig.fir 286649:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.RocketConfig.fir 286650:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.RocketConfig.fir 286645:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.RocketConfig.fir 286652:4]
      inflight_1 <= 160'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.RocketConfig.fir 286652:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.RocketConfig.fir 286925:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 286654:4]
      inflight_sizes_1 <= 640'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 286654:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.RocketConfig.fir 286933:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286689:4]
      d_first_counter_2 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 286689:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 286699:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 286700:6]
        d_first_counter_2 <= 1'h0;
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.RocketConfig.fir 286934:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.RocketConfig.fir 286934:4]
    end else if (d_first_done) begin // @[Monitor.scala 819:47 chipyard.TestHarness.RocketConfig.fir 286958:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.RocketConfig.fir 286959:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.RocketConfig.fir 286952:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285279:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285280:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285298:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285299:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285305:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285306:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285313:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285314:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285320:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285321:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285328:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285329:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285337:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285338:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285345:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285346:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285377:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285378:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285396:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285397:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285403:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285404:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285411:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285412:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285418:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285419:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285426:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285427:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285434:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285435:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285443:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285444:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285451:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285452:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285474:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285475:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285492:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285493:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285499:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285500:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285506:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285507:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285514:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285515:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285522:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285523:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285530:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285531:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285565:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285566:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285572:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285573:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285579:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285580:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285587:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285588:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285595:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285596:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285630:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285631:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285637:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285638:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285644:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285645:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285652:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285653:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285662:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285663:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285694:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285695:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285701:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285702:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285708:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285709:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285716:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285717:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285724:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285725:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285756:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285757:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285763:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285764:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285770:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285771:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285778:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285779:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285786:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285787:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285818:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285819:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285825:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285826:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285832:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285833:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285840:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285841:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285848:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285849:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285856:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 285857:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285867:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285868:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285888:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285889:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285896:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285897:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285930:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285931:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285937:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285938:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285945:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285946:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285988:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285989:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285995:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 285996:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286003:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286004:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286047:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_214 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286048:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286082:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_216 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286083:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286118:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_218 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286119:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286214:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286215:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286222:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286223:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286230:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286231:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286238:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286239:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286246:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286247:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286295:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286296:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286311:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286312:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286319:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286320:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286480:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286481:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286540:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286541:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286551:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286552:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_220 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286559:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286560:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286573:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286574:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286581:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286582:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286600:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286601:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286612:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286613:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286640:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286641:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286862:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286863:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286883:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 286884:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286947:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 286948:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[7:0];
  _RAND_10 = {5{`RANDOM}};
  inflight = _RAND_10[159:0];
  _RAND_11 = {20{`RANDOM}};
  inflight_opcodes = _RAND_11[639:0];
  _RAND_12 = {20{`RANDOM}};
  inflight_sizes = _RAND_12[639:0];
  _RAND_13 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  watchdog = _RAND_15[31:0];
  _RAND_16 = {5{`RANDOM}};
  inflight_1 = _RAND_16[159:0];
  _RAND_17 = {20{`RANDOM}};
  inflight_sizes_1 = _RAND_17[639:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  watchdog_1 = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLRAM_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 286962:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 286963:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 286964:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  input  [1:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  input  [7:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  output [1:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  output [7:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
  output [63:0] auto_in_d_bits_data // @[chipyard.TestHarness.RocketConfig.fir 286965:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire [1:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire [7:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire [1:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire [7:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
  wire [8:0] mem_RW0_addr; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_en; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_clk; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_wmode; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_wdata_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_wdata_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_wdata_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_wdata_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_wdata_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_wdata_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_wdata_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_wdata_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_rdata_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_rdata_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_rdata_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_rdata_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_rdata_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_rdata_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_rdata_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire [7:0] mem_RW0_rdata_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_wmask_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_wmask_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_wmask_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_wmask_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_wmask_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_wmask_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_wmask_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  wire  mem_RW0_wmask_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
  reg  r_full; // @[SRAM.scala 134:30 chipyard.TestHarness.RocketConfig.fir 287011:4]
  reg [1:0] r_size; // @[SRAM.scala 137:26 chipyard.TestHarness.RocketConfig.fir 287014:4]
  reg [7:0] r_source; // @[SRAM.scala 138:26 chipyard.TestHarness.RocketConfig.fir 287015:4]
  reg  r_read; // @[SRAM.scala 139:26 chipyard.TestHarness.RocketConfig.fir 287016:4]
  reg  REG; // @[SRAM.scala 321:58 chipyard.TestHarness.RocketConfig.fir 287536:4]
  reg [7:0] r_1; // @[Reg.scala 15:16 chipyard.TestHarness.RocketConfig.fir 287538:4]
  wire [7:0] r_raw_data_1 = REG ? mem_RW0_rdata_1 : r_1; // @[package.scala 79:42 chipyard.TestHarness.RocketConfig.fir 287549:4]
  reg [7:0] r_0; // @[Reg.scala 15:16 chipyard.TestHarness.RocketConfig.fir 287538:4]
  wire [7:0] r_raw_data_0 = REG ? mem_RW0_rdata_0 : r_0; // @[package.scala 79:42 chipyard.TestHarness.RocketConfig.fir 287549:4]
  reg [7:0] r_3; // @[Reg.scala 15:16 chipyard.TestHarness.RocketConfig.fir 287538:4]
  wire [7:0] r_raw_data_3 = REG ? mem_RW0_rdata_3 : r_3; // @[package.scala 79:42 chipyard.TestHarness.RocketConfig.fir 287549:4]
  reg [7:0] r_2; // @[Reg.scala 15:16 chipyard.TestHarness.RocketConfig.fir 287538:4]
  wire [7:0] r_raw_data_2 = REG ? mem_RW0_rdata_2 : r_2; // @[package.scala 79:42 chipyard.TestHarness.RocketConfig.fir 287549:4]
  wire [31:0] r_corrected_lo = {r_raw_data_3,r_raw_data_2,r_raw_data_1,r_raw_data_0}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 287079:4]
  reg [7:0] r_5; // @[Reg.scala 15:16 chipyard.TestHarness.RocketConfig.fir 287538:4]
  wire [7:0] r_raw_data_5 = REG ? mem_RW0_rdata_5 : r_5; // @[package.scala 79:42 chipyard.TestHarness.RocketConfig.fir 287549:4]
  reg [7:0] r_4; // @[Reg.scala 15:16 chipyard.TestHarness.RocketConfig.fir 287538:4]
  wire [7:0] r_raw_data_4 = REG ? mem_RW0_rdata_4 : r_4; // @[package.scala 79:42 chipyard.TestHarness.RocketConfig.fir 287549:4]
  reg [7:0] r_7; // @[Reg.scala 15:16 chipyard.TestHarness.RocketConfig.fir 287538:4]
  wire [7:0] r_raw_data_7 = REG ? mem_RW0_rdata_7 : r_7; // @[package.scala 79:42 chipyard.TestHarness.RocketConfig.fir 287549:4]
  reg [7:0] r_6; // @[Reg.scala 15:16 chipyard.TestHarness.RocketConfig.fir 287538:4]
  wire [7:0] r_raw_data_6 = REG ? mem_RW0_rdata_6 : r_6; // @[package.scala 79:42 chipyard.TestHarness.RocketConfig.fir 287549:4]
  wire [31:0] r_corrected_hi = {r_raw_data_7,r_raw_data_6,r_raw_data_5,r_raw_data_4}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 287082:4]
  wire  _bundleIn_0_a_ready_T_2 = ~r_full; // @[SRAM.scala 243:41 chipyard.TestHarness.RocketConfig.fir 287262:4]
  wire  in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.RocketConfig.fir 287263:4]
  wire  a_read = auto_in_a_bits_opcode == 3'h4; // @[SRAM.scala 251:35 chipyard.TestHarness.RocketConfig.fir 287271:4]
  wire  _GEN_22 = auto_in_d_ready ? 1'h0 : r_full; // @[SRAM.scala 273:20 chipyard.TestHarness.RocketConfig.fir 287300:4 SRAM.scala 273:29 chipyard.TestHarness.RocketConfig.fir 287301:6 SRAM.scala 134:30 chipyard.TestHarness.RocketConfig.fir 287011:4]
  wire  _T_18 = in_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 287303:4]
  wire  _T_19 = ~a_read; // @[SRAM.scala 287:13 chipyard.TestHarness.RocketConfig.fir 287317:6]
  wire  _GEN_24 = _T_18 | _GEN_22; // @[SRAM.scala 274:24 chipyard.TestHarness.RocketConfig.fir 287304:4 SRAM.scala 275:18 chipyard.TestHarness.RocketConfig.fir 287305:6]
  wire  a_lanes_lo_lo_lo = |auto_in_a_bits_mask[0]; // @[SRAM.scala 303:95 chipyard.TestHarness.RocketConfig.fir 287441:4]
  wire  a_lanes_lo_lo_hi = |auto_in_a_bits_mask[1]; // @[SRAM.scala 303:95 chipyard.TestHarness.RocketConfig.fir 287443:4]
  wire  a_lanes_lo_hi_lo = |auto_in_a_bits_mask[2]; // @[SRAM.scala 303:95 chipyard.TestHarness.RocketConfig.fir 287445:4]
  wire  a_lanes_lo_hi_hi = |auto_in_a_bits_mask[3]; // @[SRAM.scala 303:95 chipyard.TestHarness.RocketConfig.fir 287447:4]
  wire  a_lanes_hi_lo_lo = |auto_in_a_bits_mask[4]; // @[SRAM.scala 303:95 chipyard.TestHarness.RocketConfig.fir 287449:4]
  wire  a_lanes_hi_lo_hi = |auto_in_a_bits_mask[5]; // @[SRAM.scala 303:95 chipyard.TestHarness.RocketConfig.fir 287451:4]
  wire  a_lanes_hi_hi_lo = |auto_in_a_bits_mask[6]; // @[SRAM.scala 303:95 chipyard.TestHarness.RocketConfig.fir 287453:4]
  wire  a_lanes_hi_hi_hi = |auto_in_a_bits_mask[7]; // @[SRAM.scala 303:95 chipyard.TestHarness.RocketConfig.fir 287455:4]
  wire [7:0] a_lanes = {a_lanes_hi_hi_hi,a_lanes_hi_hi_lo,a_lanes_hi_lo_hi,a_lanes_hi_lo_lo,a_lanes_lo_hi_hi,
    a_lanes_lo_hi_lo,a_lanes_lo_lo_hi,a_lanes_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 287462:4]
  wire  wen = _T_18 & _T_19; // @[SRAM.scala 309:52 chipyard.TestHarness.RocketConfig.fir 287470:4]
  wire  _ren_T = ~wen; // @[SRAM.scala 310:15 chipyard.TestHarness.RocketConfig.fir 287473:4]
  wire  ren = _ren_T & _T_18; // @[SRAM.scala 310:20 chipyard.TestHarness.RocketConfig.fir 287475:4]
  wire  index_lo_lo_lo = auto_in_a_bits_address[3]; // @[SRAM.scala 320:60 chipyard.TestHarness.RocketConfig.fir 287494:4]
  wire  index_lo_lo_hi = auto_in_a_bits_address[4]; // @[SRAM.scala 320:60 chipyard.TestHarness.RocketConfig.fir 287495:4]
  wire  index_lo_hi_lo = auto_in_a_bits_address[5]; // @[SRAM.scala 320:60 chipyard.TestHarness.RocketConfig.fir 287496:4]
  wire  index_lo_hi_hi = auto_in_a_bits_address[6]; // @[SRAM.scala 320:60 chipyard.TestHarness.RocketConfig.fir 287497:4]
  wire  index_hi_lo_lo = auto_in_a_bits_address[7]; // @[SRAM.scala 320:60 chipyard.TestHarness.RocketConfig.fir 287498:4]
  wire  index_hi_lo_hi = auto_in_a_bits_address[8]; // @[SRAM.scala 320:60 chipyard.TestHarness.RocketConfig.fir 287499:4]
  wire  index_hi_hi_lo = auto_in_a_bits_address[9]; // @[SRAM.scala 320:60 chipyard.TestHarness.RocketConfig.fir 287500:4]
  wire  index_hi_hi_hi_lo = auto_in_a_bits_address[10]; // @[SRAM.scala 320:60 chipyard.TestHarness.RocketConfig.fir 287501:4]
  wire  index_hi_hi_hi_hi = auto_in_a_bits_address[11]; // @[SRAM.scala 320:60 chipyard.TestHarness.RocketConfig.fir 287502:4]
  wire [3:0] index_lo = {index_lo_hi_hi,index_lo_hi_lo,index_lo_lo_hi,index_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 287522:4]
  wire [4:0] index_hi = {index_hi_hi_hi_hi,index_hi_hi_hi_lo,index_hi_hi_lo,index_hi_lo_hi,index_hi_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 287526:4]
  TLMonitor_54_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 286972:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source)
  );
  mem_inTestHarness mem ( // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.RocketConfig.fir 286996:4]
    .RW0_addr(mem_RW0_addr),
    .RW0_en(mem_RW0_en),
    .RW0_clk(mem_RW0_clk),
    .RW0_wmode(mem_RW0_wmode),
    .RW0_wdata_0(mem_RW0_wdata_0),
    .RW0_wdata_1(mem_RW0_wdata_1),
    .RW0_wdata_2(mem_RW0_wdata_2),
    .RW0_wdata_3(mem_RW0_wdata_3),
    .RW0_wdata_4(mem_RW0_wdata_4),
    .RW0_wdata_5(mem_RW0_wdata_5),
    .RW0_wdata_6(mem_RW0_wdata_6),
    .RW0_wdata_7(mem_RW0_wdata_7),
    .RW0_rdata_0(mem_RW0_rdata_0),
    .RW0_rdata_1(mem_RW0_rdata_1),
    .RW0_rdata_2(mem_RW0_rdata_2),
    .RW0_rdata_3(mem_RW0_rdata_3),
    .RW0_rdata_4(mem_RW0_rdata_4),
    .RW0_rdata_5(mem_RW0_rdata_5),
    .RW0_rdata_6(mem_RW0_rdata_6),
    .RW0_rdata_7(mem_RW0_rdata_7),
    .RW0_wmask_0(mem_RW0_wmask_0),
    .RW0_wmask_1(mem_RW0_wmask_1),
    .RW0_wmask_2(mem_RW0_wmask_2),
    .RW0_wmask_3(mem_RW0_wmask_3),
    .RW0_wmask_4(mem_RW0_wmask_4),
    .RW0_wmask_5(mem_RW0_wmask_5),
    .RW0_wmask_6(mem_RW0_wmask_6),
    .RW0_wmask_7(mem_RW0_wmask_7)
  );
  assign auto_in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.RocketConfig.fir 287263:4]
  assign auto_in_d_valid = r_full; // @[SRAM.scala 240:65 chipyard.TestHarness.RocketConfig.fir 287242:4]
  assign auto_in_d_bits_opcode = {{2'd0}, r_read}; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 SRAM.scala 209:23 chipyard.TestHarness.RocketConfig.fir 287190:4]
  assign auto_in_d_bits_size = r_size; // @[SRAM.scala 211:29 chipyard.TestHarness.RocketConfig.fir 287192:4]
  assign auto_in_d_bits_source = r_source; // @[SRAM.scala 212:29 chipyard.TestHarness.RocketConfig.fir 287194:4]
  assign auto_in_d_bits_data = {r_corrected_hi,r_corrected_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 287090:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 286973:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 286974:4]
  assign monitor_io_in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.RocketConfig.fir 287263:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 286995:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 286995:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 286995:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 286995:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 286995:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 286995:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 286995:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 286995:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 286995:4]
  assign monitor_io_in_d_valid = r_full; // @[SRAM.scala 240:65 chipyard.TestHarness.RocketConfig.fir 287242:4]
  assign monitor_io_in_d_bits_opcode = {{2'd0}, r_read}; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 286970:4 SRAM.scala 209:23 chipyard.TestHarness.RocketConfig.fir 287190:4]
  assign monitor_io_in_d_bits_size = r_size; // @[SRAM.scala 211:29 chipyard.TestHarness.RocketConfig.fir 287192:4]
  assign monitor_io_in_d_bits_source = r_source; // @[SRAM.scala 212:29 chipyard.TestHarness.RocketConfig.fir 287194:4]
  assign mem_RW0_wdata_0 = auto_in_a_bits_data[7:0]; // @[SRAM.scala 291:67 chipyard.TestHarness.RocketConfig.fir 287322:4]
  assign mem_RW0_wdata_1 = auto_in_a_bits_data[15:8]; // @[SRAM.scala 291:67 chipyard.TestHarness.RocketConfig.fir 287323:4]
  assign mem_RW0_wdata_2 = auto_in_a_bits_data[23:16]; // @[SRAM.scala 291:67 chipyard.TestHarness.RocketConfig.fir 287324:4]
  assign mem_RW0_wdata_3 = auto_in_a_bits_data[31:24]; // @[SRAM.scala 291:67 chipyard.TestHarness.RocketConfig.fir 287325:4]
  assign mem_RW0_wdata_4 = auto_in_a_bits_data[39:32]; // @[SRAM.scala 291:67 chipyard.TestHarness.RocketConfig.fir 287326:4]
  assign mem_RW0_wdata_5 = auto_in_a_bits_data[47:40]; // @[SRAM.scala 291:67 chipyard.TestHarness.RocketConfig.fir 287327:4]
  assign mem_RW0_wdata_6 = auto_in_a_bits_data[55:48]; // @[SRAM.scala 291:67 chipyard.TestHarness.RocketConfig.fir 287328:4]
  assign mem_RW0_wdata_7 = auto_in_a_bits_data[63:56]; // @[SRAM.scala 291:67 chipyard.TestHarness.RocketConfig.fir 287329:4]
  assign mem_RW0_wmask_0 = a_lanes[0]; // @[SRAM.scala 322:46 chipyard.TestHarness.RocketConfig.fir 287559:6]
  assign mem_RW0_wmask_1 = a_lanes[1]; // @[SRAM.scala 322:46 chipyard.TestHarness.RocketConfig.fir 287560:6]
  assign mem_RW0_wmask_2 = a_lanes[2]; // @[SRAM.scala 322:46 chipyard.TestHarness.RocketConfig.fir 287561:6]
  assign mem_RW0_wmask_3 = a_lanes[3]; // @[SRAM.scala 322:46 chipyard.TestHarness.RocketConfig.fir 287562:6]
  assign mem_RW0_wmask_4 = a_lanes[4]; // @[SRAM.scala 322:46 chipyard.TestHarness.RocketConfig.fir 287563:6]
  assign mem_RW0_wmask_5 = a_lanes[5]; // @[SRAM.scala 322:46 chipyard.TestHarness.RocketConfig.fir 287564:6]
  assign mem_RW0_wmask_6 = a_lanes[6]; // @[SRAM.scala 322:46 chipyard.TestHarness.RocketConfig.fir 287565:6]
  assign mem_RW0_wmask_7 = a_lanes[7]; // @[SRAM.scala 322:46 chipyard.TestHarness.RocketConfig.fir 287566:6]
  assign mem_RW0_wmode = _T_18 & _T_19; // @[SRAM.scala 309:52 chipyard.TestHarness.RocketConfig.fir 287470:4]
  assign mem_RW0_clk = clock;
  assign mem_RW0_en = ren | wen;
  assign mem_RW0_addr = {index_hi,index_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 287527:4]
  always @(posedge clock) begin
    if (reset) begin // @[SRAM.scala 134:30 chipyard.TestHarness.RocketConfig.fir 287011:4]
      r_full <= 1'h0; // @[SRAM.scala 134:30 chipyard.TestHarness.RocketConfig.fir 287011:4]
    end else begin
      r_full <= _GEN_24;
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.RocketConfig.fir 287304:4]
      r_size <= auto_in_a_bits_size; // @[SRAM.scala 279:18 chipyard.TestHarness.RocketConfig.fir 287309:6]
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.RocketConfig.fir 287304:4]
      r_source <= auto_in_a_bits_source; // @[SRAM.scala 280:18 chipyard.TestHarness.RocketConfig.fir 287310:6]
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.RocketConfig.fir 287304:4]
      r_read <= a_read; // @[SRAM.scala 281:18 chipyard.TestHarness.RocketConfig.fir 287311:6]
    end
    REG <= _ren_T & _T_18; // @[SRAM.scala 310:20 chipyard.TestHarness.RocketConfig.fir 287475:4]
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.RocketConfig.fir 287539:4]
      r_1 <= mem_RW0_rdata_1; // @[Reg.scala 16:23 chipyard.TestHarness.RocketConfig.fir 287541:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.RocketConfig.fir 287539:4]
      r_0 <= mem_RW0_rdata_0; // @[Reg.scala 16:23 chipyard.TestHarness.RocketConfig.fir 287540:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.RocketConfig.fir 287539:4]
      r_3 <= mem_RW0_rdata_3; // @[Reg.scala 16:23 chipyard.TestHarness.RocketConfig.fir 287543:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.RocketConfig.fir 287539:4]
      r_2 <= mem_RW0_rdata_2; // @[Reg.scala 16:23 chipyard.TestHarness.RocketConfig.fir 287542:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.RocketConfig.fir 287539:4]
      r_5 <= mem_RW0_rdata_5; // @[Reg.scala 16:23 chipyard.TestHarness.RocketConfig.fir 287545:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.RocketConfig.fir 287539:4]
      r_4 <= mem_RW0_rdata_4; // @[Reg.scala 16:23 chipyard.TestHarness.RocketConfig.fir 287544:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.RocketConfig.fir 287539:4]
      r_7 <= mem_RW0_rdata_7; // @[Reg.scala 16:23 chipyard.TestHarness.RocketConfig.fir 287547:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.RocketConfig.fir 287539:4]
      r_6 <= mem_RW0_rdata_6; // @[Reg.scala 16:23 chipyard.TestHarness.RocketConfig.fir 287546:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_size = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  r_source = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  r_read = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  r_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  r_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  r_2 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  r_5 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  r_4 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  r_7 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  r_6 = _RAND_12[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar_10_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 287603:2]
  output        auto_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [2:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [3:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [2:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [3:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [2:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [3:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [2:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [3:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input         auto_out_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 287606:4]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 287611:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 287615:4]
  assign auto_in_d_valid = auto_out_d_valid; // @[ReadyValidCancel.scala 21:38 chipyard.TestHarness.RocketConfig.fir 288027:4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 287611:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 287615:4]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 287611:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 287615:4]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 287611:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 287615:4]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Xbar.scala 228:69 chipyard.TestHarness.RocketConfig.fir 287726:4]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Xbar.scala 323:53 chipyard.TestHarness.RocketConfig.fir 287788:4]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 287611:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 287615:4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 287611:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 287615:4]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 287611:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 287615:4]
  assign auto_out_a_valid = auto_in_a_valid; // @[ReadyValidCancel.scala 21:38 chipyard.TestHarness.RocketConfig.fir 288052:4]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 287613:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 287616:4]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 287613:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 287616:4]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 287613:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 287616:4]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55 chipyard.TestHarness.RocketConfig.fir 287680:4]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 287613:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 287616:4]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 287613:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 287616:4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 287613:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 287616:4]
  assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 287613:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 287616:4]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 287613:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 287616:4]
endmodule
module TLMonitor_55_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 288129:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 288130:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 288131:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input  [1:0]  io_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input  [7:0]  io_in_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input  [1:0]  io_in_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input  [7:0]  io_in_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input         io_in_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 288132:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [159:0] _RAND_13;
  reg [639:0] _RAND_14;
  reg [639:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [159:0] _RAND_19;
  reg [639:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 289623:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 289930:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.RocketConfig.fir 288149:6]
  wire [5:0] _is_aligned_mask_T_1 = 6'h7 << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 288155:6]
  wire [2:0] is_aligned_mask = ~_is_aligned_mask_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 288157:6]
  wire [28:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.RocketConfig.fir 288158:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.RocketConfig.fir 288158:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.RocketConfig.fir 288159:6]
  wire [2:0] _mask_sizeOH_T = {{1'd0}, io_in_a_bits_size}; // @[Misc.scala 201:34 chipyard.TestHarness.RocketConfig.fir 288160:6]
  wire [1:0] mask_sizeOH_shiftAmount = _mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.RocketConfig.fir 288161:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.RocketConfig.fir 288162:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.RocketConfig.fir 288164:6]
  wire  _mask_T = io_in_a_bits_size >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.RocketConfig.fir 288165:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 288166:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 288167:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 288168:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288170:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288171:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288173:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288174:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 288175:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 288176:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 288177:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288178:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288179:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288180:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288181:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288182:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288183:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288184:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288185:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288186:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288187:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288188:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288189:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 288190:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 288191:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 288192:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288193:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288194:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288195:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288196:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288197:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288198:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288199:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288200:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288201:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288202:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288203:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288204:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288205:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288206:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288207:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288208:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288209:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288210:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288211:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288212:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288213:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 288214:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 288215:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 288216:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 288223:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.RocketConfig.fir 288246:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 288262:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 288263:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 288265:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 288266:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288272:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288297:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288298:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288305:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288306:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288312:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288313:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.RocketConfig.fir 288318:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288320:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288321:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.RocketConfig.fir 288326:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.RocketConfig.fir 288327:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288329:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288330:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.RocketConfig.fir 288335:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288337:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288338:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.RocketConfig.fir 288344:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.RocketConfig.fir 288424:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288426:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288427:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.RocketConfig.fir 288450:6]
  wire  _T_175 = _T_37 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288484:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288485:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.RocketConfig.fir 288504:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288506:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288507:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.RocketConfig.fir 288512:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288514:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288515:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.RocketConfig.fir 288529:6]
  wire  _T_218 = _source_ok_T_4 & _T_37; // @[Monitor.scala 115:71 chipyard.TestHarness.RocketConfig.fir 288555:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288557:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288558:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.RocketConfig.fir 288594:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.RocketConfig.fir 288650:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.RocketConfig.fir 288651:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.RocketConfig.fir 288652:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288654:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288655:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.RocketConfig.fir 288661:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.RocketConfig.fir 288706:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288708:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288709:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.RocketConfig.fir 288723:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.RocketConfig.fir 288768:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288770:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288771:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.RocketConfig.fir 288785:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.RocketConfig.fir 288830:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288832:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288833:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.RocketConfig.fir 288857:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288859:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288860:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.RocketConfig.fir 288871:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.RocketConfig.fir 288877:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288880:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288881:8]
  wire  _T_405 = io_in_d_bits_size >= 2'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.RocketConfig.fir 288886:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288888:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288889:8]
  wire  _T_409 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.RocketConfig.fir 288894:8]
  wire  _T_411 = _T_409 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288896:8]
  wire  _T_412 = ~_T_411; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288897:8]
  wire  _T_413 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.RocketConfig.fir 288902:8]
  wire  _T_415 = _T_413 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288904:8]
  wire  _T_416 = ~_T_415; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288905:8]
  wire  _T_417 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.RocketConfig.fir 288910:8]
  wire  _T_419 = _T_417 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288912:8]
  wire  _T_420 = ~_T_419; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288913:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.RocketConfig.fir 288919:6]
  wire  _T_432 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.RocketConfig.fir 288943:8]
  wire  _T_434 = _T_432 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288945:8]
  wire  _T_435 = ~_T_434; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288946:8]
  wire  _T_436 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.RocketConfig.fir 288951:8]
  wire  _T_438 = _T_436 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288953:8]
  wire  _T_439 = ~_T_438; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288954:8]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.RocketConfig.fir 288977:6]
  wire  _T_469 = _T_417 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.RocketConfig.fir 289018:8]
  wire  _T_471 = _T_469 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289020:8]
  wire  _T_472 = ~_T_471; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289021:8]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.RocketConfig.fir 289036:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.RocketConfig.fir 289071:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.RocketConfig.fir 289107:6]
  wire  a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 289173:4]
  reg  a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289182:4]
  wire  a_first_counter1 = a_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 289184:4]
  wire  a_first = ~a_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 289185:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.RocketConfig.fir 289196:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.RocketConfig.fir 289197:4]
  reg [1:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.RocketConfig.fir 289198:4]
  reg [7:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.RocketConfig.fir 289199:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.RocketConfig.fir 289200:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.RocketConfig.fir 289201:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.RocketConfig.fir 289202:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.RocketConfig.fir 289204:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289206:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289207:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.RocketConfig.fir 289212:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289214:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289215:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.RocketConfig.fir 289220:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289222:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289223:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.RocketConfig.fir 289228:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289230:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289231:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.RocketConfig.fir 289236:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289238:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289239:6]
  wire  _T_565 = a_first_done & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.RocketConfig.fir 289246:4]
  wire  d_first_done = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 289254:4]
  reg  d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289262:4]
  wire  d_first_counter1 = d_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 289264:4]
  wire  d_first = ~d_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 289265:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.RocketConfig.fir 289276:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.RocketConfig.fir 289277:4]
  reg [1:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.RocketConfig.fir 289278:4]
  reg [7:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.RocketConfig.fir 289279:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.RocketConfig.fir 289280:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.RocketConfig.fir 289281:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.RocketConfig.fir 289282:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.RocketConfig.fir 289283:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.RocketConfig.fir 289285:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289287:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289288:6]
  wire  _T_572 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.RocketConfig.fir 289293:6]
  wire  _T_574 = _T_572 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289295:6]
  wire  _T_575 = ~_T_574; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289296:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.RocketConfig.fir 289301:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289303:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289304:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.RocketConfig.fir 289309:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289311:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289312:6]
  wire  _T_584 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.RocketConfig.fir 289317:6]
  wire  _T_586 = _T_584 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289319:6]
  wire  _T_587 = ~_T_586; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289320:6]
  wire  _T_588 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.RocketConfig.fir 289325:6]
  wire  _T_590 = _T_588 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289327:6]
  wire  _T_591 = ~_T_590; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289328:6]
  wire  _T_593 = d_first_done & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.RocketConfig.fir 289335:4]
  reg [159:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 289344:4]
  reg [639:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 289345:4]
  reg [639:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 289346:4]
  reg  a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289356:4]
  wire  a_first_counter1_1 = a_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 289358:4]
  wire  a_first_1 = ~a_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 289359:4]
  reg  d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289378:4]
  wire  d_first_counter1_1 = d_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 289380:4]
  wire  d_first_1 = ~d_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 289381:4]
  wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.RocketConfig.fir 289402:4]
  wire [10:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.RocketConfig.fir 289402:4]
  wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.RocketConfig.fir 289403:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.RocketConfig.fir 289407:4]
  wire [639:0] _GEN_73 = {{624'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.RocketConfig.fir 289408:4]
  wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.RocketConfig.fir 289408:4]
  wire [639:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[639:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.RocketConfig.fir 289409:4]
  wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.RocketConfig.fir 289414:4]
  wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.RocketConfig.fir 289419:4]
  wire [639:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[639:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.RocketConfig.fir 289420:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.RocketConfig.fir 289444:4]
  wire [255:0] _a_set_wo_ready_T = 256'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.RocketConfig.fir 289447:6]
  wire [255:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.RocketConfig.fir 289446:4 Monitor.scala 649:22 chipyard.TestHarness.RocketConfig.fir 289448:6 chipyard.TestHarness.RocketConfig.fir 289395:4]
  wire  _T_597 = a_first_done & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.RocketConfig.fir 289451:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.RocketConfig.fir 289456:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.RocketConfig.fir 289457:6]
  wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.RocketConfig.fir 289459:6]
  wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.RocketConfig.fir 289460:6]
  wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.RocketConfig.fir 289462:6]
  wire [10:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.RocketConfig.fir 289462:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 289453:4 Monitor.scala 654:28 chipyard.TestHarness.RocketConfig.fir 289458:6 chipyard.TestHarness.RocketConfig.fir 289441:4]
  wire [2050:0] _GEN_79 = {{2047'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.RocketConfig.fir 289463:6]
  wire [2050:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.RocketConfig.fir 289463:6]
  wire [2:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 3'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 289453:4 Monitor.scala 655:28 chipyard.TestHarness.RocketConfig.fir 289461:6 chipyard.TestHarness.RocketConfig.fir 289443:4]
  wire [2049:0] _GEN_81 = {{2047'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.RocketConfig.fir 289466:6]
  wire [2049:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.RocketConfig.fir 289466:6]
  wire [159:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.RocketConfig.fir 289468:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.RocketConfig.fir 289470:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289472:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289473:6]
  wire [255:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 289453:4 Monitor.scala 653:28 chipyard.TestHarness.RocketConfig.fir 289455:6 chipyard.TestHarness.RocketConfig.fir 289393:4]
  wire [2050:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 2051'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 289453:4 Monitor.scala 656:28 chipyard.TestHarness.RocketConfig.fir 289464:6 chipyard.TestHarness.RocketConfig.fir 289397:4]
  wire [2049:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 2050'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 289453:4 Monitor.scala 657:28 chipyard.TestHarness.RocketConfig.fir 289467:6 chipyard.TestHarness.RocketConfig.fir 289399:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.RocketConfig.fir 289488:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.RocketConfig.fir 289490:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.RocketConfig.fir 289491:4]
  wire [255:0] _d_clr_wo_ready_T = 256'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.RocketConfig.fir 289493:6]
  wire [255:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.RocketConfig.fir 289492:4 Monitor.scala 672:22 chipyard.TestHarness.RocketConfig.fir 289494:6 chipyard.TestHarness.RocketConfig.fir 289482:4]
  wire  _T_610 = d_first_done & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.RocketConfig.fir 289497:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.RocketConfig.fir 289500:4]
  wire [2062:0] _GEN_83 = {{2047'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.RocketConfig.fir 289509:6]
  wire [2062:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.RocketConfig.fir 289509:6]
  wire [255:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 289501:4 Monitor.scala 676:21 chipyard.TestHarness.RocketConfig.fir 289503:6 chipyard.TestHarness.RocketConfig.fir 289480:4]
  wire [2062:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 289501:4 Monitor.scala 677:21 chipyard.TestHarness.RocketConfig.fir 289510:6 chipyard.TestHarness.RocketConfig.fir 289484:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.RocketConfig.fir 289526:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.RocketConfig.fir 289527:6]
  wire [159:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.RocketConfig.fir 289528:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.RocketConfig.fir 289530:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289532:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289533:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 289539:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 289540:8 Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 289540:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 289540:8 Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 289540:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 289540:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.RocketConfig.fir 289541:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289543:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289544:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.RocketConfig.fir 289549:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289551:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289552:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 289400:4 Monitor.scala 634:21 chipyard.TestHarness.RocketConfig.fir 289410:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 289560:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 289562:8 Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 289562:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 289562:8 Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 289562:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 289562:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.RocketConfig.fir 289563:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289565:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289566:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 289411:4 Monitor.scala 638:19 chipyard.TestHarness.RocketConfig.fir 289421:4]
  wire [3:0] _GEN_86 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.RocketConfig.fir 289571:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.RocketConfig.fir 289571:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289573:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289574:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.RocketConfig.fir 289582:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.RocketConfig.fir 289583:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.RocketConfig.fir 289585:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.RocketConfig.fir 289587:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.RocketConfig.fir 289589:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.RocketConfig.fir 289590:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289592:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289593:6]
  wire [159:0] a_set_wo_ready = _GEN_15[159:0]; // @[chipyard.TestHarness.RocketConfig.fir 289394:4]
  wire [159:0] d_clr_wo_ready = _GEN_21[159:0]; // @[chipyard.TestHarness.RocketConfig.fir 289481:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.RocketConfig.fir 289599:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.RocketConfig.fir 289600:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.RocketConfig.fir 289601:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.RocketConfig.fir 289602:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289604:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289605:4]
  wire [159:0] a_set = _GEN_16[159:0]; // @[chipyard.TestHarness.RocketConfig.fir 289392:4]
  wire [159:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.RocketConfig.fir 289610:4]
  wire [159:0] d_clr = _GEN_22[159:0]; // @[chipyard.TestHarness.RocketConfig.fir 289479:4]
  wire [159:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.RocketConfig.fir 289611:4]
  wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.RocketConfig.fir 289612:4]
  wire [639:0] a_opcodes_set = _GEN_19[639:0]; // @[chipyard.TestHarness.RocketConfig.fir 289396:4]
  wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.RocketConfig.fir 289614:4]
  wire [639:0] d_opcodes_clr = _GEN_23[639:0]; // @[chipyard.TestHarness.RocketConfig.fir 289483:4]
  wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.RocketConfig.fir 289615:4]
  wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.RocketConfig.fir 289616:4]
  wire [639:0] a_sizes_set = _GEN_20[639:0]; // @[chipyard.TestHarness.RocketConfig.fir 289398:4]
  wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.RocketConfig.fir 289618:4]
  wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.RocketConfig.fir 289620:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 289622:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.RocketConfig.fir 289625:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.RocketConfig.fir 289626:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.RocketConfig.fir 289627:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.RocketConfig.fir 289628:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.RocketConfig.fir 289629:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.RocketConfig.fir 289630:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289632:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289633:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.RocketConfig.fir 289639:4]
  wire  _T_676 = a_first_done | d_first_done; // @[Monitor.scala 712:27 chipyard.TestHarness.RocketConfig.fir 289643:4]
  reg [159:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.RocketConfig.fir 289647:4]
  reg [639:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 289649:4]
  reg  d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289684:4]
  wire  d_first_counter1_2 = d_first_counter_2 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 289686:4]
  wire  d_first_2 = ~d_first_counter_2; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 289687:4]
  wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.RocketConfig.fir 289720:4]
  wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.RocketConfig.fir 289725:4]
  wire [639:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[639:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.RocketConfig.fir 289726:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.RocketConfig.fir 289804:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.RocketConfig.fir 289806:4]
  wire  _T_698 = d_first_done & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.RocketConfig.fir 289812:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.RocketConfig.fir 289814:4]
  wire [255:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.RocketConfig.fir 289815:4 Monitor.scala 784:21 chipyard.TestHarness.RocketConfig.fir 289817:6 chipyard.TestHarness.RocketConfig.fir 289796:4]
  wire [2062:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.RocketConfig.fir 289815:4 Monitor.scala 785:21 chipyard.TestHarness.RocketConfig.fir 289824:6 chipyard.TestHarness.RocketConfig.fir 289800:4]
  wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.RocketConfig.fir 289850:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289854:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289855:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 289708:4 Monitor.scala 747:21 chipyard.TestHarness.RocketConfig.fir 289727:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.RocketConfig.fir 289873:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289875:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289876:8]
  wire [159:0] d_clr_1 = _GEN_67[159:0]; // @[chipyard.TestHarness.RocketConfig.fir 289795:4]
  wire [159:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.RocketConfig.fir 289918:4]
  wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.RocketConfig.fir 289919:4]
  wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0]; // @[chipyard.TestHarness.RocketConfig.fir 289799:4]
  wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.RocketConfig.fir 289922:4]
  wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.RocketConfig.fir 289927:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.RocketConfig.fir 289929:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.RocketConfig.fir 289932:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.RocketConfig.fir 289933:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.RocketConfig.fir 289934:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.RocketConfig.fir 289935:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.RocketConfig.fir 289936:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.RocketConfig.fir 289937:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289939:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289940:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.RocketConfig.fir 289946:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288274:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288372:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288469:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288560:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288625:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288689:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288751:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288813:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288883:10]
  wire  _GEN_208 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288925:10]
  wire  _GEN_222 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288983:10]
  wire  _GEN_236 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289042:10]
  wire  _GEN_244 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289077:10]
  wire  _GEN_252 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289113:10]
  wire  _GEN_260 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289546:10]
  wire  _GEN_265 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289568:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 289623:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 289930:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289182:4]
      a_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289182:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 289192:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 289193:6]
        a_first_counter <= 1'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 289247:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.RocketConfig.fir 289248:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 289247:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.RocketConfig.fir 289249:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 289247:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.RocketConfig.fir 289250:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 289247:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.RocketConfig.fir 289251:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 289247:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.RocketConfig.fir 289252:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289262:4]
      d_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289262:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 289272:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 289273:6]
        d_first_counter <= 1'h0;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 289336:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.RocketConfig.fir 289337:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 289336:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.RocketConfig.fir 289338:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 289336:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.RocketConfig.fir 289339:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 289336:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.RocketConfig.fir 289340:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 289336:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.RocketConfig.fir 289341:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 289336:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.RocketConfig.fir 289342:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 289344:4]
      inflight <= 160'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 289344:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.RocketConfig.fir 289613:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 289345:4]
      inflight_opcodes <= 640'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 289345:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.RocketConfig.fir 289617:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 289346:4]
      inflight_sizes <= 640'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 289346:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.RocketConfig.fir 289621:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289356:4]
      a_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289356:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 289366:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 289367:6]
        a_first_counter_1 <= 1'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289378:4]
      d_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289378:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 289388:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 289389:6]
        d_first_counter_1 <= 1'h0;
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 289622:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 289622:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.RocketConfig.fir 289644:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.RocketConfig.fir 289645:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.RocketConfig.fir 289640:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.RocketConfig.fir 289647:4]
      inflight_1 <= 160'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.RocketConfig.fir 289647:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.RocketConfig.fir 289920:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 289649:4]
      inflight_sizes_1 <= 640'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 289649:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.RocketConfig.fir 289928:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289684:4]
      d_first_counter_2 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 289684:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 289694:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 289695:6]
        d_first_counter_2 <= 1'h0;
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.RocketConfig.fir 289929:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.RocketConfig.fir 289929:4]
    end else if (d_first_done) begin // @[Monitor.scala 819:47 chipyard.TestHarness.RocketConfig.fir 289953:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.RocketConfig.fir 289954:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.RocketConfig.fir 289947:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288274:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288275:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288293:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288294:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288300:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288301:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288308:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288309:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288315:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288316:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288323:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288324:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288332:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288333:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288340:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288341:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288372:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288373:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288391:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288392:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288398:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288399:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288406:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288407:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288413:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288414:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288421:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288422:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288429:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288430:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288438:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288439:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288446:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288447:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288469:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288470:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288487:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288488:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288494:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288495:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288501:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288502:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288509:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288510:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288517:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288518:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288525:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288526:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288560:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288561:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288567:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288568:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288574:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288575:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288582:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288583:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288590:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288591:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288625:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288626:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288632:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288633:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288639:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288640:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288647:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288648:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288657:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288658:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288689:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288690:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288696:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288697:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288703:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288704:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288711:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288712:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288719:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288720:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288751:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288752:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288758:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288759:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288765:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288766:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288773:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288774:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288781:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288782:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288813:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288814:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288820:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288821:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288827:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288828:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288835:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288836:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288843:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288844:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288851:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 288852:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288862:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288863:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288883:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288884:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288891:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288892:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288899:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288900:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288907:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288908:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288915:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288916:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288925:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288926:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288932:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288933:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288940:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288941:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288948:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288949:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288956:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288957:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288964:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288965:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288973:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288974:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288983:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288984:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288990:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288991:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288998:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 288999:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289006:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289007:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289014:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289015:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289023:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289024:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289032:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289033:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289042:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289043:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289050:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289051:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289058:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289059:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289067:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289068:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289077:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289078:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289085:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289086:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289094:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289095:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289103:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289104:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289113:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289114:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289121:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289122:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289129:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289130:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289138:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289139:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289209:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289210:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289217:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289218:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289225:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289226:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289233:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289234:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289241:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289242:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289290:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289291:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289298:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289299:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289306:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289307:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289314:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289315:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289322:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289323:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289330:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289331:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289475:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289476:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289535:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289536:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289546:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289547:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289554:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289555:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289568:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289569:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289576:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289577:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289595:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289596:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289607:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289608:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289635:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289636:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289857:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289858:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289878:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 289879:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289942:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 289943:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {5{`RANDOM}};
  inflight = _RAND_13[159:0];
  _RAND_14 = {20{`RANDOM}};
  inflight_opcodes = _RAND_14[639:0];
  _RAND_15 = {20{`RANDOM}};
  inflight_sizes = _RAND_15[639:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {5{`RANDOM}};
  inflight_1 = _RAND_19[159:0];
  _RAND_20 = {20{`RANDOM}};
  inflight_sizes_1 = _RAND_20[639:0];
  _RAND_21 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  watchdog_1 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_40_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 289957:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 289958:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 289959:4]
  output        io_enq_ready, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  input         io_enq_valid, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  input  [2:0]  io_enq_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  input  [1:0]  io_enq_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  input  [7:0]  io_enq_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  input  [28:0] io_enq_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  input  [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  input         io_deq_ready, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  output        io_deq_valid, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  output [1:0]  io_deq_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  output [7:0]  io_deq_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  output [28:0] io_deq_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  output [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 289960:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  reg [1:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  reg [7:0] ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [7:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [7:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  reg [28:0] ram_address [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [28:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [28:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 289963:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 289964:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 289965:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.RocketConfig.fir 289966:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.RocketConfig.fir 289967:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.RocketConfig.fir 289968:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.RocketConfig.fir 289969:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 289970:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 289973:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 289988:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 289994:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.RocketConfig.fir 289997:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.RocketConfig.fir 290003:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.RocketConfig.fir 290001:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290013:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290012:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290011:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290010:4]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290009:4]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290008:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290007:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290006:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 289962:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 289963:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 289963:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.RocketConfig.fir 289976:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 289989:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 289964:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 289964:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.RocketConfig.fir 289991:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 289995:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 289965:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 289965:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.RocketConfig.fir 289998:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.RocketConfig.fir 289999:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[28:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_41_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 290021:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 290022:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 290023:4]
  output        io_enq_ready, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  input         io_enq_valid, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  input  [1:0]  io_enq_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  input  [7:0]  io_enq_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  input         io_deq_ready, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  output        io_deq_valid, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  output [1:0]  io_deq_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  output [1:0]  io_deq_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  output [7:0]  io_deq_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  output        io_deq_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  output        io_deq_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 290024:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  reg [1:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  reg [7:0] ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire [7:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire [7:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  reg  ram_sink [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 290027:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 290028:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 290029:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.RocketConfig.fir 290030:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.RocketConfig.fir 290031:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.RocketConfig.fir 290032:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.RocketConfig.fir 290033:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 290034:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 290037:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 290052:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 290058:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.RocketConfig.fir 290061:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  assign ram_param_MPORT_data = 2'h0;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_addr = value_1;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  assign ram_sink_MPORT_data = 1'h0;
  assign ram_sink_MPORT_addr = value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  assign ram_denied_MPORT_data = 1'h0;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.RocketConfig.fir 290067:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.RocketConfig.fir 290065:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290077:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290076:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290075:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290074:4]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290073:4]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290072:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290071:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 290070:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 290026:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 290027:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 290027:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.RocketConfig.fir 290040:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 290053:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 290028:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 290028:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.RocketConfig.fir 290055:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 290059:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 290029:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 290029:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.RocketConfig.fir 290062:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.RocketConfig.fir 290063:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_20_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 290085:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 290086:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 290087:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [1:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [7:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [1:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [7:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [1:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [7:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [1:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [7:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
  input  [63:0] auto_out_d_bits_data // @[chipyard.TestHarness.RocketConfig.fir 290088:4]
);
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire [1:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire [7:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire [1:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire [7:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [1:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [28:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire  bundleOut_0_a_q_io_enq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [1:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [28:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire  bundleOut_0_a_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire [1:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire [7:0] bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire [7:0] bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire  bundleIn_0_d_q_io_deq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
  TLMonitor_55_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 290095:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_40_inTestHarness bundleOut_0_a_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290122:4]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
  );
  Queue_41_inTestHarness bundleIn_0_d_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 290136:4]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Decoupled.scala 299:17 chipyard.TestHarness.RocketConfig.fir 290134:4]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 290135:4]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 290135:4]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 290135:4]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 290135:4]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 290135:4]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 290135:4]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 290135:4]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 290135:4]
  assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 290135:4]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 Decoupled.scala 299:17 chipyard.TestHarness.RocketConfig.fir 290148:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 290096:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 290097:4]
  assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Decoupled.scala 299:17 chipyard.TestHarness.RocketConfig.fir 290134:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 290149:4]
  assign bundleOut_0_a_q_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 290123:4]
  assign bundleOut_0_a_q_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 290124:4]
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 290120:4]
  assign bundleIn_0_d_q_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 290137:4]
  assign bundleIn_0_d_q_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 290138:4]
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 290120:4]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 290120:4]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 290120:4]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 290120:4]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 290118:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 290120:4]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 290093:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 290121:4]
endmodule
module TLMonitor_56_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 290185:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 290186:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 290187:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input  [2:0]  io_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input  [3:0]  io_in_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input  [2:0]  io_in_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input  [3:0]  io_in_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input         io_in_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 290188:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 291679:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 291986:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 4'h9; // @[Parameters.scala 57:20 chipyard.TestHarness.RocketConfig.fir 290205:6]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 290211:6]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 290213:6]
  wire [28:0] _GEN_71 = {{23'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.RocketConfig.fir 290214:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.RocketConfig.fir 290214:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.RocketConfig.fir 290215:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.RocketConfig.fir 290217:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.RocketConfig.fir 290218:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.RocketConfig.fir 290220:6]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21 chipyard.TestHarness.RocketConfig.fir 290221:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 290222:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 290223:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 290224:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290226:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290227:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290229:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290230:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 290231:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 290232:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 290233:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290234:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290235:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290236:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290237:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290238:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290239:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290240:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290241:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290242:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290243:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290244:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290245:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 290246:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 290247:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 290248:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290249:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290250:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290251:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290252:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290253:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290254:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290255:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290256:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290257:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290258:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290259:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290260:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290261:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290262:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290263:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290264:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290265:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290266:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290267:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290268:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290269:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 290270:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 290271:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 290272:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 290279:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.RocketConfig.fir 290302:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 290318:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 290319:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 290321:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 290322:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290328:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290353:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290354:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290361:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290362:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290368:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290369:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.RocketConfig.fir 290374:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290376:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290377:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.RocketConfig.fir 290382:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.RocketConfig.fir 290383:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290385:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290386:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.RocketConfig.fir 290391:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290393:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290394:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.RocketConfig.fir 290400:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.RocketConfig.fir 290480:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290482:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290483:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.RocketConfig.fir 290506:6]
  wire  _T_164 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.RocketConfig.fir 290529:8]
  wire  _T_172 = _T_164 & _T_37; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 290537:8]
  wire  _T_175 = _T_172 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290540:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290541:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.RocketConfig.fir 290560:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290562:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290563:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.RocketConfig.fir 290568:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290570:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290571:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.RocketConfig.fir 290585:6]
  wire  _T_218 = _source_ok_T_4 & _T_172; // @[Monitor.scala 115:71 chipyard.TestHarness.RocketConfig.fir 290611:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290613:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290614:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.RocketConfig.fir 290650:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.RocketConfig.fir 290706:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.RocketConfig.fir 290707:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.RocketConfig.fir 290708:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290710:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290711:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.RocketConfig.fir 290717:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.RocketConfig.fir 290762:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290764:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290765:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.RocketConfig.fir 290779:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.RocketConfig.fir 290824:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290826:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290827:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.RocketConfig.fir 290841:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.RocketConfig.fir 290886:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290888:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290889:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.RocketConfig.fir 290913:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290915:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290916:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 4'h9; // @[Parameters.scala 57:20 chipyard.TestHarness.RocketConfig.fir 290927:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.RocketConfig.fir 290933:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290936:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290937:8]
  wire  _T_405 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.RocketConfig.fir 290942:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290944:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290945:8]
  wire  _T_409 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.RocketConfig.fir 290950:8]
  wire  _T_411 = _T_409 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290952:8]
  wire  _T_412 = ~_T_411; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290953:8]
  wire  _T_413 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.RocketConfig.fir 290958:8]
  wire  _T_415 = _T_413 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290960:8]
  wire  _T_416 = ~_T_415; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290961:8]
  wire  _T_417 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.RocketConfig.fir 290966:8]
  wire  _T_419 = _T_417 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290968:8]
  wire  _T_420 = ~_T_419; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290969:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.RocketConfig.fir 290975:6]
  wire  _T_432 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.RocketConfig.fir 290999:8]
  wire  _T_434 = _T_432 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291001:8]
  wire  _T_435 = ~_T_434; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291002:8]
  wire  _T_436 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.RocketConfig.fir 291007:8]
  wire  _T_438 = _T_436 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291009:8]
  wire  _T_439 = ~_T_438; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291010:8]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.RocketConfig.fir 291033:6]
  wire  _T_469 = _T_417 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.RocketConfig.fir 291074:8]
  wire  _T_471 = _T_469 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291076:8]
  wire  _T_472 = ~_T_471; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291077:8]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.RocketConfig.fir 291092:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.RocketConfig.fir 291127:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.RocketConfig.fir 291163:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 291229:4]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.RocketConfig.fir 291234:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.RocketConfig.fir 291236:4]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291238:4]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 291240:4]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 291241:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.RocketConfig.fir 291252:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.RocketConfig.fir 291253:4]
  reg [2:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.RocketConfig.fir 291254:4]
  reg [3:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.RocketConfig.fir 291255:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.RocketConfig.fir 291256:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.RocketConfig.fir 291257:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.RocketConfig.fir 291258:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.RocketConfig.fir 291260:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291262:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291263:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.RocketConfig.fir 291268:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291270:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291271:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.RocketConfig.fir 291276:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291278:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291279:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.RocketConfig.fir 291284:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291286:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291287:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.RocketConfig.fir 291292:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291294:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291295:6]
  wire  _T_565 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.RocketConfig.fir 291302:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 291310:4]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 291312:4]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 291314:4]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.RocketConfig.fir 291315:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.RocketConfig.fir 291316:4]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291318:4]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 291320:4]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 291321:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.RocketConfig.fir 291332:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.RocketConfig.fir 291333:4]
  reg [2:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.RocketConfig.fir 291334:4]
  reg [3:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.RocketConfig.fir 291335:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.RocketConfig.fir 291336:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.RocketConfig.fir 291337:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.RocketConfig.fir 291338:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.RocketConfig.fir 291339:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.RocketConfig.fir 291341:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291343:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291344:6]
  wire  _T_572 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.RocketConfig.fir 291349:6]
  wire  _T_574 = _T_572 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291351:6]
  wire  _T_575 = ~_T_574; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291352:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.RocketConfig.fir 291357:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291359:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291360:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.RocketConfig.fir 291365:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291367:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291368:6]
  wire  _T_584 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.RocketConfig.fir 291373:6]
  wire  _T_586 = _T_584 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291375:6]
  wire  _T_587 = ~_T_586; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291376:6]
  wire  _T_588 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.RocketConfig.fir 291381:6]
  wire  _T_590 = _T_588 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291383:6]
  wire  _T_591 = ~_T_590; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291384:6]
  wire  _T_593 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.RocketConfig.fir 291391:4]
  reg [9:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 291400:4]
  reg [39:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 291401:4]
  reg [39:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 291402:4]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291412:4]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 291414:4]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 291415:4]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291434:4]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 291436:4]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 291437:4]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.RocketConfig.fir 291458:4]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.RocketConfig.fir 291458:4]
  wire [39:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.RocketConfig.fir 291459:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.RocketConfig.fir 291463:4]
  wire [39:0] _GEN_73 = {{24'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.RocketConfig.fir 291464:4]
  wire [39:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.RocketConfig.fir 291464:4]
  wire [39:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[39:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.RocketConfig.fir 291465:4]
  wire [39:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.RocketConfig.fir 291470:4]
  wire [39:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.RocketConfig.fir 291475:4]
  wire [39:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[39:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.RocketConfig.fir 291476:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.RocketConfig.fir 291500:4]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.RocketConfig.fir 291503:6]
  wire [15:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.RocketConfig.fir 291502:4 Monitor.scala 649:22 chipyard.TestHarness.RocketConfig.fir 291504:6 chipyard.TestHarness.RocketConfig.fir 291451:4]
  wire  _T_597 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.RocketConfig.fir 291507:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.RocketConfig.fir 291512:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.RocketConfig.fir 291513:6]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.RocketConfig.fir 291515:6]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.RocketConfig.fir 291516:6]
  wire [5:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.RocketConfig.fir 291518:6]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.RocketConfig.fir 291518:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 291509:4 Monitor.scala 654:28 chipyard.TestHarness.RocketConfig.fir 291514:6 chipyard.TestHarness.RocketConfig.fir 291497:4]
  wire [130:0] _GEN_79 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.RocketConfig.fir 291519:6]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.RocketConfig.fir 291519:6]
  wire [3:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 291509:4 Monitor.scala 655:28 chipyard.TestHarness.RocketConfig.fir 291517:6 chipyard.TestHarness.RocketConfig.fir 291499:4]
  wire [130:0] _GEN_81 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.RocketConfig.fir 291522:6]
  wire [130:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.RocketConfig.fir 291522:6]
  wire [9:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.RocketConfig.fir 291524:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.RocketConfig.fir 291526:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291528:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291529:6]
  wire [15:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 291509:4 Monitor.scala 653:28 chipyard.TestHarness.RocketConfig.fir 291511:6 chipyard.TestHarness.RocketConfig.fir 291449:4]
  wire [130:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 291509:4 Monitor.scala 656:28 chipyard.TestHarness.RocketConfig.fir 291520:6 chipyard.TestHarness.RocketConfig.fir 291453:4]
  wire [130:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 291509:4 Monitor.scala 657:28 chipyard.TestHarness.RocketConfig.fir 291523:6 chipyard.TestHarness.RocketConfig.fir 291455:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.RocketConfig.fir 291544:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.RocketConfig.fir 291546:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.RocketConfig.fir 291547:4]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.RocketConfig.fir 291549:6]
  wire [15:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.RocketConfig.fir 291548:4 Monitor.scala 672:22 chipyard.TestHarness.RocketConfig.fir 291550:6 chipyard.TestHarness.RocketConfig.fir 291538:4]
  wire  _T_610 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.RocketConfig.fir 291553:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.RocketConfig.fir 291556:4]
  wire [142:0] _GEN_83 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.RocketConfig.fir 291565:6]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.RocketConfig.fir 291565:6]
  wire [15:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 291557:4 Monitor.scala 676:21 chipyard.TestHarness.RocketConfig.fir 291559:6 chipyard.TestHarness.RocketConfig.fir 291536:4]
  wire [142:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 291557:4 Monitor.scala 677:21 chipyard.TestHarness.RocketConfig.fir 291566:6 chipyard.TestHarness.RocketConfig.fir 291540:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.RocketConfig.fir 291582:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.RocketConfig.fir 291583:6]
  wire [9:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.RocketConfig.fir 291584:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.RocketConfig.fir 291586:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291588:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291589:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 291595:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 291596:8 Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 291596:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 291596:8 Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 291596:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 291596:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.RocketConfig.fir 291597:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291599:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291600:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.RocketConfig.fir 291605:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291607:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291608:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 291456:4 Monitor.scala 634:21 chipyard.TestHarness.RocketConfig.fir 291466:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 291616:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 291618:8 Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 291618:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 291618:8 Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 291618:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 291618:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.RocketConfig.fir 291619:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291621:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291622:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 291467:4 Monitor.scala 638:19 chipyard.TestHarness.RocketConfig.fir 291477:4]
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.RocketConfig.fir 291627:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.RocketConfig.fir 291627:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291629:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291630:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.RocketConfig.fir 291638:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.RocketConfig.fir 291639:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.RocketConfig.fir 291641:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.RocketConfig.fir 291643:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.RocketConfig.fir 291645:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.RocketConfig.fir 291646:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291648:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291649:6]
  wire [9:0] a_set_wo_ready = _GEN_15[9:0]; // @[chipyard.TestHarness.RocketConfig.fir 291450:4]
  wire [9:0] d_clr_wo_ready = _GEN_21[9:0]; // @[chipyard.TestHarness.RocketConfig.fir 291537:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.RocketConfig.fir 291655:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.RocketConfig.fir 291656:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.RocketConfig.fir 291657:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.RocketConfig.fir 291658:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291660:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291661:4]
  wire [9:0] a_set = _GEN_16[9:0]; // @[chipyard.TestHarness.RocketConfig.fir 291448:4]
  wire [9:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.RocketConfig.fir 291666:4]
  wire [9:0] d_clr = _GEN_22[9:0]; // @[chipyard.TestHarness.RocketConfig.fir 291535:4]
  wire [9:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.RocketConfig.fir 291667:4]
  wire [9:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.RocketConfig.fir 291668:4]
  wire [39:0] a_opcodes_set = _GEN_19[39:0]; // @[chipyard.TestHarness.RocketConfig.fir 291452:4]
  wire [39:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.RocketConfig.fir 291670:4]
  wire [39:0] d_opcodes_clr = _GEN_23[39:0]; // @[chipyard.TestHarness.RocketConfig.fir 291539:4]
  wire [39:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.RocketConfig.fir 291671:4]
  wire [39:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.RocketConfig.fir 291672:4]
  wire [39:0] a_sizes_set = _GEN_20[39:0]; // @[chipyard.TestHarness.RocketConfig.fir 291454:4]
  wire [39:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.RocketConfig.fir 291674:4]
  wire [39:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.RocketConfig.fir 291676:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 291678:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.RocketConfig.fir 291681:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.RocketConfig.fir 291682:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.RocketConfig.fir 291683:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.RocketConfig.fir 291684:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.RocketConfig.fir 291685:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.RocketConfig.fir 291686:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291688:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291689:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.RocketConfig.fir 291695:4]
  wire  _T_676 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.RocketConfig.fir 291699:4]
  reg [9:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.RocketConfig.fir 291703:4]
  reg [39:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 291705:4]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291740:4]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 291742:4]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 291743:4]
  wire [39:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.RocketConfig.fir 291776:4]
  wire [39:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.RocketConfig.fir 291781:4]
  wire [39:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[39:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.RocketConfig.fir 291782:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.RocketConfig.fir 291860:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.RocketConfig.fir 291862:4]
  wire  _T_698 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.RocketConfig.fir 291868:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.RocketConfig.fir 291870:4]
  wire [15:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.RocketConfig.fir 291871:4 Monitor.scala 784:21 chipyard.TestHarness.RocketConfig.fir 291873:6 chipyard.TestHarness.RocketConfig.fir 291852:4]
  wire [142:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.RocketConfig.fir 291871:4 Monitor.scala 785:21 chipyard.TestHarness.RocketConfig.fir 291880:6 chipyard.TestHarness.RocketConfig.fir 291856:4]
  wire [9:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.RocketConfig.fir 291906:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291910:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291911:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 291764:4 Monitor.scala 747:21 chipyard.TestHarness.RocketConfig.fir 291783:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.RocketConfig.fir 291929:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291931:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291932:8]
  wire [9:0] d_clr_1 = _GEN_67[9:0]; // @[chipyard.TestHarness.RocketConfig.fir 291851:4]
  wire [9:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.RocketConfig.fir 291974:4]
  wire [9:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.RocketConfig.fir 291975:4]
  wire [39:0] d_opcodes_clr_1 = _GEN_68[39:0]; // @[chipyard.TestHarness.RocketConfig.fir 291855:4]
  wire [39:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.RocketConfig.fir 291978:4]
  wire [39:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.RocketConfig.fir 291983:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.RocketConfig.fir 291985:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.RocketConfig.fir 291988:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.RocketConfig.fir 291989:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.RocketConfig.fir 291990:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.RocketConfig.fir 291991:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.RocketConfig.fir 291992:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.RocketConfig.fir 291993:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291995:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291996:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.RocketConfig.fir 292002:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290330:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290428:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290525:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290616:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290681:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290745:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290807:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290869:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290939:10]
  wire  _GEN_208 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290981:10]
  wire  _GEN_222 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291039:10]
  wire  _GEN_236 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291098:10]
  wire  _GEN_244 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291133:10]
  wire  _GEN_252 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291169:10]
  wire  _GEN_260 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291602:10]
  wire  _GEN_265 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291624:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 291679:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 291986:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291238:4]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291238:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 291248:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 291249:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 291237:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 291303:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.RocketConfig.fir 291304:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 291303:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.RocketConfig.fir 291305:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 291303:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.RocketConfig.fir 291306:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 291303:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.RocketConfig.fir 291307:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 291303:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.RocketConfig.fir 291308:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291318:4]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291318:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 291328:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 291329:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 291317:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 291392:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.RocketConfig.fir 291393:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 291392:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.RocketConfig.fir 291394:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 291392:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.RocketConfig.fir 291395:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 291392:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.RocketConfig.fir 291396:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 291392:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.RocketConfig.fir 291397:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 291392:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.RocketConfig.fir 291398:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 291400:4]
      inflight <= 10'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 291400:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.RocketConfig.fir 291669:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 291401:4]
      inflight_opcodes <= 40'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 291401:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.RocketConfig.fir 291673:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 291402:4]
      inflight_sizes <= 40'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 291402:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.RocketConfig.fir 291677:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291412:4]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291412:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 291422:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 291423:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 291237:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291434:4]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291434:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 291444:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 291445:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 291317:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 291678:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 291678:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.RocketConfig.fir 291700:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.RocketConfig.fir 291701:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.RocketConfig.fir 291696:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.RocketConfig.fir 291703:4]
      inflight_1 <= 10'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.RocketConfig.fir 291703:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.RocketConfig.fir 291976:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 291705:4]
      inflight_sizes_1 <= 40'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 291705:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.RocketConfig.fir 291984:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291740:4]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 291740:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 291750:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 291751:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 291317:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.RocketConfig.fir 291985:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.RocketConfig.fir 291985:4]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47 chipyard.TestHarness.RocketConfig.fir 292009:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.RocketConfig.fir 292010:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.RocketConfig.fir 292003:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290330:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290331:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290349:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290350:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290356:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290357:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290364:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290365:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290371:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290372:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290379:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290380:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290388:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290389:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290396:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290397:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290428:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290429:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290447:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290448:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290454:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290455:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290462:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290463:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290469:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290470:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290477:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290478:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290485:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290486:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290494:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290495:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290502:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290503:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290525:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290526:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290543:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290544:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290550:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290551:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290557:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290558:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290565:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290566:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290573:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290574:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290581:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290582:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290616:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290617:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290623:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290624:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290630:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290631:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290638:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290639:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290646:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290647:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290681:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290682:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290688:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290689:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290695:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290696:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290703:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290704:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290713:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290714:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290745:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290746:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290752:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290753:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290759:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290760:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290767:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290768:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290775:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290776:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290807:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290808:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290814:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290815:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290821:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290822:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290829:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290830:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290837:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290838:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290869:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290870:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290876:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290877:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290883:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290884:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290891:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290892:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290899:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290900:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290907:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 290908:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290918:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290919:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290939:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290940:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290947:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290948:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290955:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290956:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290963:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290964:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290971:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290972:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290981:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290982:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290988:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290989:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290996:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 290997:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291004:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291005:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291012:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291013:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291020:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291021:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291029:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291030:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291039:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291040:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291046:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291047:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291054:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291055:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291062:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291063:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291070:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291071:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291079:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291080:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291088:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291089:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291098:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291099:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291106:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291107:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291114:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291115:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291123:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291124:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291133:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291134:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291141:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291142:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291150:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291151:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291159:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291160:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291169:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291170:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291177:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291178:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291185:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291186:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291194:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291195:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291265:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291266:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291273:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291274:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291281:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291282:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291289:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291290:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291297:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291298:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291346:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291347:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291354:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291355:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291362:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291363:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291370:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291371:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291378:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291379:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291386:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291387:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291531:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291532:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291591:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291592:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291602:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291603:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291610:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291611:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291624:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291625:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291632:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291633:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291651:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291652:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291663:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291664:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291691:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291692:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291913:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291914:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291934:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 291935:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291998:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 291999:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[9:0];
  _RAND_14 = {2{`RANDOM}};
  inflight_opcodes = _RAND_14[39:0];
  _RAND_15 = {2{`RANDOM}};
  inflight_sizes = _RAND_15[39:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_1 = _RAND_19[9:0];
  _RAND_20 = {2{`RANDOM}};
  inflight_sizes_1 = _RAND_20[39:0];
  _RAND_21 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  watchdog_1 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater_7_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 292013:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 292014:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 292015:4]
  input         io_repeat, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  output        io_full, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  output        io_enq_ready, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  input         io_enq_valid, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  input  [2:0]  io_enq_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  input  [2:0]  io_enq_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  input  [3:0]  io_enq_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  input  [28:0] io_enq_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  input  [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  input         io_deq_ready, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  output        io_deq_valid, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  output [2:0]  io_deq_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  output [3:0]  io_deq_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  output [28:0] io_deq_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  output [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 292016:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21 chipyard.TestHarness.RocketConfig.fir 292018:4]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18 chipyard.TestHarness.RocketConfig.fir 292019:4]
  reg [2:0] saved_param; // @[Repeater.scala 20:18 chipyard.TestHarness.RocketConfig.fir 292019:4]
  reg [2:0] saved_size; // @[Repeater.scala 20:18 chipyard.TestHarness.RocketConfig.fir 292019:4]
  reg [3:0] saved_source; // @[Repeater.scala 20:18 chipyard.TestHarness.RocketConfig.fir 292019:4]
  reg [28:0] saved_address; // @[Repeater.scala 20:18 chipyard.TestHarness.RocketConfig.fir 292019:4]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18 chipyard.TestHarness.RocketConfig.fir 292019:4]
  reg  saved_corrupt; // @[Repeater.scala 20:18 chipyard.TestHarness.RocketConfig.fir 292019:4]
  wire  _io_enq_ready_T = ~full; // @[Repeater.scala 24:35 chipyard.TestHarness.RocketConfig.fir 292022:4]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 292035:4]
  wire  _T_1 = _T & io_repeat; // @[Repeater.scala 28:23 chipyard.TestHarness.RocketConfig.fir 292036:4]
  wire  _GEN_0 = _T_1 | full; // @[Repeater.scala 28:38 chipyard.TestHarness.RocketConfig.fir 292037:4 Repeater.scala 28:45 chipyard.TestHarness.RocketConfig.fir 292038:6 Repeater.scala 19:21 chipyard.TestHarness.RocketConfig.fir 292018:4]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 292048:4]
  wire  _T_3 = ~io_repeat; // @[Repeater.scala 29:26 chipyard.TestHarness.RocketConfig.fir 292049:4]
  wire  _T_4 = _T_2 & _T_3; // @[Repeater.scala 29:23 chipyard.TestHarness.RocketConfig.fir 292050:4]
  assign io_full = full; // @[Repeater.scala 26:11 chipyard.TestHarness.RocketConfig.fir 292034:4]
  assign io_enq_ready = io_deq_ready & _io_enq_ready_T; // @[Repeater.scala 24:32 chipyard.TestHarness.RocketConfig.fir 292023:4]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32 chipyard.TestHarness.RocketConfig.fir 292020:4]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21 chipyard.TestHarness.RocketConfig.fir 292025:4]
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; // @[Repeater.scala 25:21 chipyard.TestHarness.RocketConfig.fir 292025:4]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21 chipyard.TestHarness.RocketConfig.fir 292025:4]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21 chipyard.TestHarness.RocketConfig.fir 292025:4]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21 chipyard.TestHarness.RocketConfig.fir 292025:4]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21 chipyard.TestHarness.RocketConfig.fir 292025:4]
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; // @[Repeater.scala 25:21 chipyard.TestHarness.RocketConfig.fir 292025:4]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21 chipyard.TestHarness.RocketConfig.fir 292018:4]
      full <= 1'h0; // @[Repeater.scala 19:21 chipyard.TestHarness.RocketConfig.fir 292018:4]
    end else if (_T_4) begin // @[Repeater.scala 29:38 chipyard.TestHarness.RocketConfig.fir 292051:4]
      full <= 1'h0; // @[Repeater.scala 29:45 chipyard.TestHarness.RocketConfig.fir 292052:6]
    end else begin
      full <= _GEN_0;
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.RocketConfig.fir 292037:4]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62 chipyard.TestHarness.RocketConfig.fir 292046:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.RocketConfig.fir 292037:4]
      saved_param <= io_enq_bits_param; // @[Repeater.scala 28:62 chipyard.TestHarness.RocketConfig.fir 292045:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.RocketConfig.fir 292037:4]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62 chipyard.TestHarness.RocketConfig.fir 292044:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.RocketConfig.fir 292037:4]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62 chipyard.TestHarness.RocketConfig.fir 292043:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.RocketConfig.fir 292037:4]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62 chipyard.TestHarness.RocketConfig.fir 292042:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.RocketConfig.fir 292037:4]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62 chipyard.TestHarness.RocketConfig.fir 292041:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.RocketConfig.fir 292037:4]
      saved_corrupt <= io_enq_bits_corrupt; // @[Repeater.scala 28:62 chipyard.TestHarness.RocketConfig.fir 292039:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  saved_address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  saved_mask = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  saved_corrupt = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter_8_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 292055:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 292056:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 292057:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [2:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [3:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [2:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [3:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [1:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [7:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [1:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [7:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input         auto_out_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 292058:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
  wire  repeater_clock; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire  repeater_reset; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [2:0] repeater_io_enq_bits_opcode; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [2:0] repeater_io_enq_bits_param; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [3:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [28:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [7:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire  repeater_io_enq_bits_corrupt; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [2:0] repeater_io_deq_bits_opcode; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [2:0] repeater_io_deq_bits_param; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [3:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [28:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire [7:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  wire  repeater_io_deq_bits_corrupt; // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
  reg [2:0] acknum; // @[Fragmenter.scala 189:29 chipyard.TestHarness.RocketConfig.fir 292092:4]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24 chipyard.TestHarness.RocketConfig.fir 292093:4]
  reg  dToggle; // @[Fragmenter.scala 191:30 chipyard.TestHarness.RocketConfig.fir 292094:4]
  wire [2:0] dFragnum = auto_out_d_bits_source[2:0]; // @[Fragmenter.scala 192:41 chipyard.TestHarness.RocketConfig.fir 292095:4]
  wire  dFirst = acknum == 3'h0; // @[Fragmenter.scala 193:29 chipyard.TestHarness.RocketConfig.fir 292096:4]
  wire  dLast = dFragnum == 3'h0; // @[Fragmenter.scala 194:30 chipyard.TestHarness.RocketConfig.fir 292097:4]
  wire [3:0] dsizeOH = 4'h1 << auto_out_d_bits_size; // @[OneHot.scala 65:12 chipyard.TestHarness.RocketConfig.fir 292099:4]
  wire [5:0] _dsizeOH1_T_1 = 6'h7 << auto_out_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 292102:4]
  wire [2:0] dsizeOH1 = ~_dsizeOH1_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 292104:4]
  wire  dHasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.RocketConfig.fir 292105:4]
  wire  ack_decrement = dHasData | dsizeOH[3]; // @[Fragmenter.scala 204:32 chipyard.TestHarness.RocketConfig.fir 292122:4]
  wire [5:0] _dFirst_size_T = {dFragnum, 3'h0}; // @[Fragmenter.scala 206:47 chipyard.TestHarness.RocketConfig.fir 292123:4]
  wire [5:0] _GEN_7 = {{3'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69 chipyard.TestHarness.RocketConfig.fir 292124:4]
  wire [5:0] dFirst_size_lo = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69 chipyard.TestHarness.RocketConfig.fir 292124:4]
  wire [6:0] _dFirst_size_T_1 = {dFirst_size_lo, 1'h0}; // @[package.scala 232:35 chipyard.TestHarness.RocketConfig.fir 292125:4]
  wire [6:0] _dFirst_size_T_2 = _dFirst_size_T_1 | 7'h1; // @[package.scala 232:40 chipyard.TestHarness.RocketConfig.fir 292126:4]
  wire [6:0] _dFirst_size_T_3 = {1'h0,dFirst_size_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 292127:4]
  wire [6:0] _dFirst_size_T_4 = ~_dFirst_size_T_3; // @[package.scala 232:53 chipyard.TestHarness.RocketConfig.fir 292128:4]
  wire [6:0] _dFirst_size_T_5 = _dFirst_size_T_2 & _dFirst_size_T_4; // @[package.scala 232:51 chipyard.TestHarness.RocketConfig.fir 292129:4]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_5[6:4]; // @[OneHot.scala 30:18 chipyard.TestHarness.RocketConfig.fir 292130:4]
  wire [3:0] dFirst_size_lo_1 = _dFirst_size_T_5[3:0]; // @[OneHot.scala 31:18 chipyard.TestHarness.RocketConfig.fir 292131:4]
  wire  dFirst_size_hi_1 = |dFirst_size_hi; // @[OneHot.scala 32:14 chipyard.TestHarness.RocketConfig.fir 292132:4]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28 chipyard.TestHarness.RocketConfig.fir 292133:4]
  wire [3:0] _dFirst_size_T_6 = _GEN_8 | dFirst_size_lo_1; // @[OneHot.scala 32:28 chipyard.TestHarness.RocketConfig.fir 292133:4]
  wire [1:0] dFirst_size_hi_2 = _dFirst_size_T_6[3:2]; // @[OneHot.scala 30:18 chipyard.TestHarness.RocketConfig.fir 292134:4]
  wire [1:0] dFirst_size_lo_2 = _dFirst_size_T_6[1:0]; // @[OneHot.scala 31:18 chipyard.TestHarness.RocketConfig.fir 292135:4]
  wire  dFirst_size_hi_3 = |dFirst_size_hi_2; // @[OneHot.scala 32:14 chipyard.TestHarness.RocketConfig.fir 292136:4]
  wire [1:0] _dFirst_size_T_7 = dFirst_size_hi_2 | dFirst_size_lo_2; // @[OneHot.scala 32:28 chipyard.TestHarness.RocketConfig.fir 292137:4]
  wire  dFirst_size_lo_3 = _dFirst_size_T_7[1]; // @[CircuitMath.scala 30:8 chipyard.TestHarness.RocketConfig.fir 292138:4]
  wire [2:0] dFirst_size = {dFirst_size_hi_1,dFirst_size_hi_3,dFirst_size_lo_3}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 292140:4]
  wire  _drop_T = ~dHasData; // @[Fragmenter.scala 222:20 chipyard.TestHarness.RocketConfig.fir 292153:4]
  wire  _drop_T_2 = ~dLast; // @[Fragmenter.scala 222:33 chipyard.TestHarness.RocketConfig.fir 292155:4]
  wire  drop = _drop_T & _drop_T_2; // @[Fragmenter.scala 222:30 chipyard.TestHarness.RocketConfig.fir 292156:4]
  wire  bundleOut_0_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35 chipyard.TestHarness.RocketConfig.fir 292157:4]
  wire  _T_7 = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 292141:4]
  wire [2:0] _GEN_9 = {{2'd0}, ack_decrement}; // @[Fragmenter.scala 209:55 chipyard.TestHarness.RocketConfig.fir 292143:6]
  wire [2:0] _acknum_T_1 = acknum - _GEN_9; // @[Fragmenter.scala 209:55 chipyard.TestHarness.RocketConfig.fir 292144:6]
  wire  _bundleIn_0_d_valid_T = ~drop; // @[Fragmenter.scala 224:39 chipyard.TestHarness.RocketConfig.fir 292159:4]
  wire  _aFrag_T = repeater_io_deq_bits_size > 3'h3; // @[Fragmenter.scala 285:31 chipyard.TestHarness.RocketConfig.fir 292192:4]
  wire [2:0] aFrag = _aFrag_T ? 3'h3 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24 chipyard.TestHarness.RocketConfig.fir 292193:4]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 292195:4]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 292197:4]
  wire [9:0] _aFragOH1_T_1 = 10'h7 << aFrag; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 292199:4]
  wire [2:0] aFragOH1 = ~_aFragOH1_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 292201:4]
  wire  aHasData = ~repeater_io_deq_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.RocketConfig.fir 292203:4]
  reg [2:0] gennum; // @[Fragmenter.scala 291:29 chipyard.TestHarness.RocketConfig.fir 292205:4]
  wire  aFirst = gennum == 3'h0; // @[Fragmenter.scala 292:29 chipyard.TestHarness.RocketConfig.fir 292206:4]
  wire [2:0] _old_gennum1_T_2 = gennum - 3'h1; // @[Fragmenter.scala 293:79 chipyard.TestHarness.RocketConfig.fir 292209:4]
  wire [2:0] old_gennum1 = aFirst ? aOrigOH1[5:3] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30 chipyard.TestHarness.RocketConfig.fir 292210:4]
  wire [2:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28 chipyard.TestHarness.RocketConfig.fir 292211:4]
  wire [2:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26 chipyard.TestHarness.RocketConfig.fir 292214:4]
  reg  aToggle_r; // @[Reg.scala 15:16 chipyard.TestHarness.RocketConfig.fir 292221:4]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:19 chipyard.TestHarness.RocketConfig.fir 292222:4 Reg.scala 16:23 chipyard.TestHarness.RocketConfig.fir 292223:6 Reg.scala 15:16 chipyard.TestHarness.RocketConfig.fir 292221:4]
  wire  bundleOut_0_a_bits_source_hi_lo = ~_GEN_5; // @[Fragmenter.scala 297:23 chipyard.TestHarness.RocketConfig.fir 292226:4]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 Fragmenter.scala 303:15 chipyard.TestHarness.RocketConfig.fir 292235:4]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 292227:4]
  wire  _repeater_io_repeat_T = ~aHasData; // @[Fragmenter.scala 302:31 chipyard.TestHarness.RocketConfig.fir 292231:4]
  wire  _repeater_io_repeat_T_1 = new_gennum != 3'h0; // @[Fragmenter.scala 302:53 chipyard.TestHarness.RocketConfig.fir 292232:4]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 3'h0}; // @[Fragmenter.scala 304:65 chipyard.TestHarness.RocketConfig.fir 292236:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90 chipyard.TestHarness.RocketConfig.fir 292237:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88 chipyard.TestHarness.RocketConfig.fir 292238:4]
  wire [5:0] _GEN_10 = {{3'd0}, aFragOH1}; // @[Fragmenter.scala 304:100 chipyard.TestHarness.RocketConfig.fir 292239:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10; // @[Fragmenter.scala 304:100 chipyard.TestHarness.RocketConfig.fir 292239:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h7; // @[Fragmenter.scala 304:111 chipyard.TestHarness.RocketConfig.fir 292240:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51 chipyard.TestHarness.RocketConfig.fir 292241:4]
  wire [28:0] _GEN_11 = {{23'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49 chipyard.TestHarness.RocketConfig.fir 292242:4]
  wire [4:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,bundleOut_0_a_bits_source_hi_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 292244:4]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17 chipyard.TestHarness.RocketConfig.fir 292248:4]
  wire  _T_11 = _T_9 | _repeater_io_repeat_T; // @[Fragmenter.scala 309:35 chipyard.TestHarness.RocketConfig.fir 292250:4]
  wire  _T_13 = _T_11 | reset; // @[Fragmenter.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292252:4]
  wire  _T_14 = ~_T_13; // @[Fragmenter.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292253:4]
  wire  _T_16 = repeater_io_deq_bits_mask == 8'hff; // @[Fragmenter.scala 312:53 chipyard.TestHarness.RocketConfig.fir 292260:4]
  wire  _T_17 = _T_9 | _T_16; // @[Fragmenter.scala 312:35 chipyard.TestHarness.RocketConfig.fir 292261:4]
  wire  _T_19 = _T_17 | reset; // @[Fragmenter.scala 312:16 chipyard.TestHarness.RocketConfig.fir 292263:4]
  wire  _T_20 = ~_T_19; // @[Fragmenter.scala 312:16 chipyard.TestHarness.RocketConfig.fir 292264:4]
  TLMonitor_56_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 292065:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Repeater_7_inTestHarness repeater ( // @[Fragmenter.scala 262:30 chipyard.TestHarness.RocketConfig.fir 292167:4]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_opcode(repeater_io_enq_bits_opcode),
    .io_enq_bits_param(repeater_io_enq_bits_param),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_opcode(repeater_io_deq_bits_opcode),
    .io_deq_bits_param(repeater_io_deq_bits_param),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 Fragmenter.scala 263:25 chipyard.TestHarness.RocketConfig.fir 292171:4]
  assign auto_in_d_valid = auto_out_d_valid & _bundleIn_0_d_valid_T; // @[Fragmenter.scala 224:36 chipyard.TestHarness.RocketConfig.fir 292160:4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32 chipyard.TestHarness.RocketConfig.fir 292165:4]
  assign auto_in_d_bits_source = auto_out_d_bits_source[7:4]; // @[Fragmenter.scala 226:47 chipyard.TestHarness.RocketConfig.fir 292163:4]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 Fragmenter.scala 303:15 chipyard.TestHarness.RocketConfig.fir 292235:4]
  assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 Fragmenter.scala 303:15 chipyard.TestHarness.RocketConfig.fir 292235:4]
  assign auto_out_a_bits_param = repeater_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 Fragmenter.scala 303:15 chipyard.TestHarness.RocketConfig.fir 292235:4]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 Fragmenter.scala 306:25 chipyard.TestHarness.RocketConfig.fir 292247:4]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 292245:4]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11; // @[Fragmenter.scala 304:49 chipyard.TestHarness.RocketConfig.fir 292242:4]
  assign auto_out_a_bits_mask = repeater_io_full ? 8'hff : auto_in_a_bits_mask; // @[Fragmenter.scala 313:31 chipyard.TestHarness.RocketConfig.fir 292269:4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 Fragmenter.scala 303:15 chipyard.TestHarness.RocketConfig.fir 292235:4]
  assign auto_out_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35 chipyard.TestHarness.RocketConfig.fir 292157:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 292066:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 292067:4]
  assign monitor_io_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 Fragmenter.scala 263:25 chipyard.TestHarness.RocketConfig.fir 292171:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign monitor_io_in_d_valid = auto_out_d_valid & _bundleIn_0_d_valid_T; // @[Fragmenter.scala 224:36 chipyard.TestHarness.RocketConfig.fir 292160:4]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign monitor_io_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32 chipyard.TestHarness.RocketConfig.fir 292165:4]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:4]; // @[Fragmenter.scala 226:47 chipyard.TestHarness.RocketConfig.fir 292163:4]
  assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  assign repeater_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 292169:4]
  assign repeater_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 292170:4]
  assign repeater_io_repeat = _repeater_io_repeat_T & _repeater_io_repeat_T_1; // @[Fragmenter.scala 302:41 chipyard.TestHarness.RocketConfig.fir 292233:4]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign repeater_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 292063:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292091:4]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 292088:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 292090:4]
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29 chipyard.TestHarness.RocketConfig.fir 292092:4]
      acknum <= 3'h0; // @[Fragmenter.scala 189:29 chipyard.TestHarness.RocketConfig.fir 292092:4]
    end else if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.RocketConfig.fir 292142:4]
      if (dFirst) begin // @[Fragmenter.scala 209:24 chipyard.TestHarness.RocketConfig.fir 292145:6]
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.RocketConfig.fir 292142:4]
      if (dFirst) begin // @[Fragmenter.scala 210:25 chipyard.TestHarness.RocketConfig.fir 292147:6]
        dOrig <= dFirst_size; // @[Fragmenter.scala 211:19 chipyard.TestHarness.RocketConfig.fir 292148:8]
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30 chipyard.TestHarness.RocketConfig.fir 292094:4]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30 chipyard.TestHarness.RocketConfig.fir 292094:4]
    end else if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.RocketConfig.fir 292142:4]
      if (dFirst) begin // @[Fragmenter.scala 210:25 chipyard.TestHarness.RocketConfig.fir 292147:6]
        dToggle <= auto_out_d_bits_source[3]; // @[Fragmenter.scala 212:21 chipyard.TestHarness.RocketConfig.fir 292150:8]
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29 chipyard.TestHarness.RocketConfig.fir 292205:4]
      gennum <= 3'h0; // @[Fragmenter.scala 291:29 chipyard.TestHarness.RocketConfig.fir 292205:4]
    end else if (_T_8) begin // @[Fragmenter.scala 300:29 chipyard.TestHarness.RocketConfig.fir 292228:4]
      gennum <= new_gennum; // @[Fragmenter.scala 300:38 chipyard.TestHarness.RocketConfig.fir 292229:6]
    end
    if (aFirst) begin // @[Reg.scala 16:19 chipyard.TestHarness.RocketConfig.fir 292222:4]
      aToggle_r <= dToggle; // @[Reg.scala 16:23 chipyard.TestHarness.RocketConfig.fir 292223:6]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:309 assert (!repeater.io.full || !aHasData)\n"
            ); // @[Fragmenter.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292255:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_14) begin
          $fatal; // @[Fragmenter.scala 309:16 chipyard.TestHarness.RocketConfig.fir 292256:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16 chipyard.TestHarness.RocketConfig.fir 292266:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_20) begin
          $fatal; // @[Fragmenter.scala 312:16 chipyard.TestHarness.RocketConfig.fir 292267:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_57_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 292307:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 292308:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 292309:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input  [3:0]  io_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input  [31:0] io_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input  [3:0]  io_in_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input         io_in_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input  [2:0]  io_in_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 292310:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 294249:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 294556:4]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 292326:6]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 292328:6]
  wire [31:0] _GEN_71 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.RocketConfig.fir 292329:6]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.RocketConfig.fir 292329:6]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24 chipyard.TestHarness.RocketConfig.fir 292330:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.RocketConfig.fir 292332:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.RocketConfig.fir 292333:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.RocketConfig.fir 292335:6]
  wire  _mask_T = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21 chipyard.TestHarness.RocketConfig.fir 292336:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 292337:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 292338:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 292339:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292341:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292342:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292344:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292345:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 292346:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 292347:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 292348:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292349:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292350:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292351:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292352:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292353:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292354:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292355:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292356:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292357:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292358:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292359:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292360:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.RocketConfig.fir 292361:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.RocketConfig.fir 292362:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.RocketConfig.fir 292363:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292364:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292365:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292366:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292367:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292368:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292369:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292370:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292371:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292372:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292373:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292374:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292375:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292376:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292377:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292378:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292379:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292380:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292381:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292382:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292383:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292384:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.RocketConfig.fir 292385:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.RocketConfig.fir 292386:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.RocketConfig.fir 292387:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.RocketConfig.fir 292394:6]
  wire [32:0] _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 292398:6]
  wire  _T_15 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.RocketConfig.fir 292410:6]
  wire  _T_17 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42 chipyard.TestHarness.RocketConfig.fir 292413:8]
  wire [32:0] _T_26 = $signed(_T_7) & -33'sh101000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 292422:8]
  wire  _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 292423:8]
  wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 292424:8]
  wire [32:0] _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 292425:8]
  wire [32:0] _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 292427:8]
  wire  _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 292428:8]
  wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 292429:8]
  wire [32:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 292430:8]
  wire [32:0] _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 292432:8]
  wire  _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 292433:8]
  wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 292434:8]
  wire [32:0] _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 292435:8]
  wire [32:0] _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 292437:8]
  wire  _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 292438:8]
  wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h2010000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 292439:8]
  wire [32:0] _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 292440:8]
  wire [32:0] _T_46 = $signed(_T_44) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 292442:8]
  wire  _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 292443:8]
  wire [31:0] _T_48 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 292444:8]
  wire [32:0] _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 292445:8]
  wire [32:0] _T_51 = $signed(_T_49) & -33'sh4000000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 292447:8]
  wire  _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 292448:8]
  wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h54000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 292449:8]
  wire [32:0] _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 292450:8]
  wire [32:0] _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 292452:8]
  wire  _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 292453:8]
  wire  _T_58 = _T_27 | _T_32; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292454:8]
  wire  _T_65 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48 chipyard.TestHarness.RocketConfig.fir 292461:8]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 292463:8]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 292464:8]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 292466:8]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 292467:8]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31 chipyard.TestHarness.RocketConfig.fir 292468:8]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49 chipyard.TestHarness.RocketConfig.fir 292469:8]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh10000000; // @[Parameters.scala 137:52 chipyard.TestHarness.RocketConfig.fir 292471:8]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.RocketConfig.fir 292472:8]
  wire  _T_77 = _T_71 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292473:8]
  wire  _T_78 = _T_65 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 292474:8]
  wire  _T_81 = _T_17 & _T_78; // @[Monitor.scala 82:72 chipyard.TestHarness.RocketConfig.fir 292477:8]
  wire  _T_83 = _T_81 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292479:8]
  wire  _T_84 = ~_T_83; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292480:8]
  wire  _T_147 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292547:8]
  wire  _T_153 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292561:8]
  wire  _T_154 = ~_T_153; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292562:8]
  wire  _T_156 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292568:8]
  wire  _T_157 = ~_T_156; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292569:8]
  wire [7:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.RocketConfig.fir 292582:8]
  wire  _T_163 = _T_162 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.RocketConfig.fir 292583:8]
  wire  _T_165 = _T_163 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292585:8]
  wire  _T_166 = ~_T_165; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292586:8]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.RocketConfig.fir 292600:6]
  wire  _T_331 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.RocketConfig.fir 292798:6]
  wire  _T_339 = _T_17 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292807:8]
  wire  _T_340 = ~_T_339; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292808:8]
  wire  _T_350 = _T_17 & _T_32; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 292822:8]
  wire  _T_352 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.RocketConfig.fir 292824:8]
  wire  _T_395 = _T_27 | _T_37; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292867:8]
  wire  _T_396 = _T_395 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292868:8]
  wire  _T_397 = _T_396 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292869:8]
  wire  _T_398 = _T_397 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292870:8]
  wire  _T_399 = _T_398 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292871:8]
  wire  _T_400 = _T_399 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292872:8]
  wire  _T_401 = _T_400 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292873:8]
  wire  _T_402 = _T_352 & _T_401; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 292874:8]
  wire  _T_404 = _T_350 | _T_402; // @[Parameters.scala 672:30 chipyard.TestHarness.RocketConfig.fir 292876:8]
  wire  _T_406 = _T_404 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292878:8]
  wire  _T_407 = ~_T_406; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292879:8]
  wire  _T_418 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.RocketConfig.fir 292906:8]
  wire  _T_420 = _T_418 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292908:8]
  wire  _T_421 = ~_T_420; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292909:8]
  wire  _T_426 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.RocketConfig.fir 292923:6]
  wire  _T_482 = _T_27 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292980:8]
  wire  _T_483 = _T_482 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292981:8]
  wire  _T_484 = _T_483 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292982:8]
  wire  _T_485 = _T_484 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292983:8]
  wire  _T_486 = _T_485 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292984:8]
  wire  _T_487 = _T_486 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 292985:8]
  wire  _T_488 = _T_352 & _T_487; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 292986:8]
  wire  _T_497 = _T_350 | _T_488; // @[Parameters.scala 672:30 chipyard.TestHarness.RocketConfig.fir 292995:8]
  wire  _T_499 = _T_17 & _T_497; // @[Monitor.scala 115:71 chipyard.TestHarness.RocketConfig.fir 292997:8]
  wire  _T_501 = _T_499 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292999:8]
  wire  _T_502 = ~_T_501; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293000:8]
  wire  _T_517 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.RocketConfig.fir 293036:6]
  wire [7:0] _T_604 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.RocketConfig.fir 293140:8]
  wire [7:0] _T_605 = io_in_a_bits_mask & _T_604; // @[Monitor.scala 127:31 chipyard.TestHarness.RocketConfig.fir 293141:8]
  wire  _T_606 = _T_605 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.RocketConfig.fir 293142:8]
  wire  _T_608 = _T_606 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293144:8]
  wire  _T_609 = ~_T_608; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293145:8]
  wire  _T_610 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.RocketConfig.fir 293151:6]
  wire  _T_618 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 92:42 chipyard.TestHarness.RocketConfig.fir 293160:8]
  wire  _T_662 = _T_58 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 293204:8]
  wire  _T_663 = _T_662 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 293205:8]
  wire  _T_664 = _T_663 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 293206:8]
  wire  _T_665 = _T_664 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 293207:8]
  wire  _T_666 = _T_665 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 293208:8]
  wire  _T_667 = _T_666 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.RocketConfig.fir 293209:8]
  wire  _T_668 = _T_618 & _T_667; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 293210:8]
  wire  _T_678 = _T_17 & _T_668; // @[Monitor.scala 131:74 chipyard.TestHarness.RocketConfig.fir 293220:8]
  wire  _T_680 = _T_678 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293222:8]
  wire  _T_681 = ~_T_680; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293223:8]
  wire  _T_696 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.RocketConfig.fir 293259:6]
  wire  _T_782 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.RocketConfig.fir 293367:6]
  wire  _T_851 = _T_352 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.RocketConfig.fir 293437:8]
  wire  _T_854 = _T_350 | _T_851; // @[Parameters.scala 672:30 chipyard.TestHarness.RocketConfig.fir 293440:8]
  wire  _T_855 = _T_17 & _T_854; // @[Monitor.scala 147:68 chipyard.TestHarness.RocketConfig.fir 293441:8]
  wire  _T_857 = _T_855 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293443:8]
  wire  _T_858 = ~_T_857; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293444:8]
  wire  _T_877 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.RocketConfig.fir 293490:6]
  wire  _T_879 = _T_877 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293492:6]
  wire  _T_880 = ~_T_879; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293493:6]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.RocketConfig.fir 293498:6]
  wire  _T_881 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.RocketConfig.fir 293503:6]
  wire  _T_883 = _source_ok_T_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293506:8]
  wire  _T_884 = ~_T_883; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293507:8]
  wire  _T_885 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.RocketConfig.fir 293512:8]
  wire  _T_887 = _T_885 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293514:8]
  wire  _T_888 = ~_T_887; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293515:8]
  wire  _T_889 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.RocketConfig.fir 293520:8]
  wire  _T_891 = _T_889 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293522:8]
  wire  _T_892 = ~_T_891; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293523:8]
  wire  _T_893 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.RocketConfig.fir 293528:8]
  wire  _T_895 = _T_893 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293530:8]
  wire  _T_896 = ~_T_895; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293531:8]
  wire  _T_897 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.RocketConfig.fir 293536:8]
  wire  _T_899 = _T_897 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293538:8]
  wire  _T_900 = ~_T_899; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293539:8]
  wire  _T_901 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.RocketConfig.fir 293545:6]
  wire  _T_912 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.RocketConfig.fir 293569:8]
  wire  _T_914 = _T_912 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293571:8]
  wire  _T_915 = ~_T_914; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293572:8]
  wire  _T_916 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.RocketConfig.fir 293577:8]
  wire  _T_918 = _T_916 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293579:8]
  wire  _T_919 = ~_T_918; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293580:8]
  wire  _T_929 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.RocketConfig.fir 293603:6]
  wire  _T_949 = _T_897 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.RocketConfig.fir 293644:8]
  wire  _T_951 = _T_949 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293646:8]
  wire  _T_952 = ~_T_951; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293647:8]
  wire  _T_958 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.RocketConfig.fir 293662:6]
  wire  _T_975 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.RocketConfig.fir 293697:6]
  wire  _T_993 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.RocketConfig.fir 293733:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 293799:4]
  wire [8:0] a_first_beats1_decode = is_aligned_mask[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.RocketConfig.fir 293804:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.RocketConfig.fir 293806:4]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 293808:4]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 293810:4]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 293811:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.RocketConfig.fir 293822:4]
  reg [3:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.RocketConfig.fir 293824:4]
  reg [31:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.RocketConfig.fir 293826:4]
  wire  _T_1022 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.RocketConfig.fir 293827:4]
  wire  _T_1023 = io_in_a_valid & _T_1022; // @[Monitor.scala 389:19 chipyard.TestHarness.RocketConfig.fir 293828:4]
  wire  _T_1024 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.RocketConfig.fir 293830:6]
  wire  _T_1026 = _T_1024 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293832:6]
  wire  _T_1027 = ~_T_1026; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293833:6]
  wire  _T_1032 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.RocketConfig.fir 293846:6]
  wire  _T_1034 = _T_1032 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293848:6]
  wire  _T_1035 = ~_T_1034; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293849:6]
  wire  _T_1040 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.RocketConfig.fir 293862:6]
  wire  _T_1042 = _T_1040 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293864:6]
  wire  _T_1043 = ~_T_1042; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293865:6]
  wire  _T_1045 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.RocketConfig.fir 293872:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 293880:4]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.RocketConfig.fir 293882:4]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.RocketConfig.fir 293884:4]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.RocketConfig.fir 293885:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.RocketConfig.fir 293886:4]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 293888:4]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 293890:4]
  wire  d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 293891:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.RocketConfig.fir 293902:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.RocketConfig.fir 293903:4]
  reg [3:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.RocketConfig.fir 293904:4]
  reg  source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.RocketConfig.fir 293905:4]
  reg [2:0] sink; // @[Monitor.scala 539:22 chipyard.TestHarness.RocketConfig.fir 293906:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.RocketConfig.fir 293907:4]
  wire  _T_1046 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.RocketConfig.fir 293908:4]
  wire  _T_1047 = io_in_d_valid & _T_1046; // @[Monitor.scala 541:19 chipyard.TestHarness.RocketConfig.fir 293909:4]
  wire  _T_1048 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.RocketConfig.fir 293911:6]
  wire  _T_1050 = _T_1048 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293913:6]
  wire  _T_1051 = ~_T_1050; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293914:6]
  wire  _T_1052 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.RocketConfig.fir 293919:6]
  wire  _T_1054 = _T_1052 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293921:6]
  wire  _T_1055 = ~_T_1054; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293922:6]
  wire  _T_1056 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.RocketConfig.fir 293927:6]
  wire  _T_1058 = _T_1056 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293929:6]
  wire  _T_1059 = ~_T_1058; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293930:6]
  wire  _T_1060 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.RocketConfig.fir 293935:6]
  wire  _T_1062 = _T_1060 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293937:6]
  wire  _T_1063 = ~_T_1062; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293938:6]
  wire  _T_1064 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.RocketConfig.fir 293943:6]
  wire  _T_1066 = _T_1064 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293945:6]
  wire  _T_1067 = ~_T_1066; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293946:6]
  wire  _T_1068 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.RocketConfig.fir 293951:6]
  wire  _T_1070 = _T_1068 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293953:6]
  wire  _T_1071 = ~_T_1070; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293954:6]
  wire  _T_1073 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.RocketConfig.fir 293961:4]
  reg  inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 293970:4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 293971:4]
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 293972:4]
  reg [8:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 293982:4]
  wire [8:0] a_first_counter1_1 = a_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 293984:4]
  wire  a_first_1 = a_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 293985:4]
  reg [8:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 294004:4]
  wire [8:0] d_first_counter1_1 = d_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 294006:4]
  wire  d_first_1 = d_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 294007:4]
  wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.RocketConfig.fir 294028:4]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.RocketConfig.fir 294028:4]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.RocketConfig.fir 294029:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.RocketConfig.fir 294033:4]
  wire [15:0] _GEN_73 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.RocketConfig.fir 294034:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.RocketConfig.fir 294034:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.RocketConfig.fir 294035:4]
  wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65 chipyard.TestHarness.RocketConfig.fir 294039:4]
  wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.RocketConfig.fir 294040:4]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.RocketConfig.fir 294044:4]
  wire [15:0] _GEN_75 = {{8'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.RocketConfig.fir 294045:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.RocketConfig.fir 294045:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.RocketConfig.fir 294046:4]
  wire  _T_1074 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.RocketConfig.fir 294070:4]
  wire [1:0] _GEN_15 = _T_1074 ? 2'h1 : 2'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.RocketConfig.fir 294072:4 Monitor.scala 649:22 chipyard.TestHarness.RocketConfig.fir 294074:6 chipyard.TestHarness.RocketConfig.fir 294021:4]
  wire  _T_1077 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.RocketConfig.fir 294077:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.RocketConfig.fir 294082:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.RocketConfig.fir 294083:6]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.RocketConfig.fir 294085:6]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.RocketConfig.fir 294086:6]
  wire [3:0] a_opcodes_set_interm = _T_1077 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 294079:4 Monitor.scala 654:28 chipyard.TestHarness.RocketConfig.fir 294084:6 chipyard.TestHarness.RocketConfig.fir 294067:4]
  wire [18:0] _a_opcodes_set_T_1 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.RocketConfig.fir 294089:6]
  wire [4:0] a_sizes_set_interm = _T_1077 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 294079:4 Monitor.scala 655:28 chipyard.TestHarness.RocketConfig.fir 294087:6 chipyard.TestHarness.RocketConfig.fir 294069:4]
  wire [19:0] _a_sizes_set_T_1 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.RocketConfig.fir 294092:6]
  wire  _T_1081 = ~inflight; // @[Monitor.scala 658:17 chipyard.TestHarness.RocketConfig.fir 294096:6]
  wire  _T_1083 = _T_1081 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 294098:6]
  wire  _T_1084 = ~_T_1083; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 294099:6]
  wire [1:0] _GEN_16 = _T_1077 ? 2'h1 : 2'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 294079:4 Monitor.scala 653:28 chipyard.TestHarness.RocketConfig.fir 294081:6 chipyard.TestHarness.RocketConfig.fir 294019:4]
  wire [18:0] _GEN_19 = _T_1077 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 294079:4 Monitor.scala 656:28 chipyard.TestHarness.RocketConfig.fir 294090:6 chipyard.TestHarness.RocketConfig.fir 294023:4]
  wire [19:0] _GEN_20 = _T_1077 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.RocketConfig.fir 294079:4 Monitor.scala 657:28 chipyard.TestHarness.RocketConfig.fir 294093:6 chipyard.TestHarness.RocketConfig.fir 294025:4]
  wire  _T_1085 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.RocketConfig.fir 294114:4]
  wire  _T_1087 = ~_T_881; // @[Monitor.scala 671:74 chipyard.TestHarness.RocketConfig.fir 294116:4]
  wire  _T_1088 = _T_1085 & _T_1087; // @[Monitor.scala 671:71 chipyard.TestHarness.RocketConfig.fir 294117:4]
  wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.RocketConfig.fir 294119:6]
  wire [1:0] _GEN_21 = _T_1088 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.RocketConfig.fir 294118:4 Monitor.scala 672:22 chipyard.TestHarness.RocketConfig.fir 294120:6 chipyard.TestHarness.RocketConfig.fir 294108:4]
  wire  _T_1090 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.RocketConfig.fir 294123:4]
  wire  _T_1093 = _T_1090 & _T_1087; // @[Monitor.scala 675:72 chipyard.TestHarness.RocketConfig.fir 294126:4]
  wire [30:0] _GEN_78 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.RocketConfig.fir 294135:6]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_78 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.RocketConfig.fir 294135:6]
  wire [30:0] _GEN_79 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74 chipyard.TestHarness.RocketConfig.fir 294142:6]
  wire [30:0] _d_sizes_clr_T_5 = _GEN_79 << _a_size_lookup_T; // @[Monitor.scala 678:74 chipyard.TestHarness.RocketConfig.fir 294142:6]
  wire [1:0] _GEN_22 = _T_1093 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 294127:4 Monitor.scala 676:21 chipyard.TestHarness.RocketConfig.fir 294129:6 chipyard.TestHarness.RocketConfig.fir 294106:4]
  wire [30:0] _GEN_23 = _T_1093 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 294127:4 Monitor.scala 677:21 chipyard.TestHarness.RocketConfig.fir 294136:6 chipyard.TestHarness.RocketConfig.fir 294110:4]
  wire [30:0] _GEN_24 = _T_1093 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.RocketConfig.fir 294127:4 Monitor.scala 678:21 chipyard.TestHarness.RocketConfig.fir 294143:6 chipyard.TestHarness.RocketConfig.fir 294112:4]
  wire  same_cycle_resp = _T_1074 & _source_ok_T_1; // @[Monitor.scala 681:88 chipyard.TestHarness.RocketConfig.fir 294153:6]
  wire  _T_1098 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.RocketConfig.fir 294154:6]
  wire  _T_1100 = _T_1098 | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.RocketConfig.fir 294156:6]
  wire  _T_1102 = _T_1100 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294158:6]
  wire  _T_1103 = ~_T_1102; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294159:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8 Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8]
  wire  _T_1104 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.RocketConfig.fir 294165:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 294166:8 Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 294166:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 294166:8 Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 294166:8]
  wire  _T_1105 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.RocketConfig.fir 294166:8]
  wire  _T_1106 = _T_1104 | _T_1105; // @[Monitor.scala 685:77 chipyard.TestHarness.RocketConfig.fir 294167:8]
  wire  _T_1108 = _T_1106 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294169:8]
  wire  _T_1109 = ~_T_1108; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294170:8]
  wire  _T_1110 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.RocketConfig.fir 294175:8]
  wire  _T_1112 = _T_1110 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294177:8]
  wire  _T_1113 = ~_T_1112; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294178:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 294026:4 Monitor.scala 634:21 chipyard.TestHarness.RocketConfig.fir 294036:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8 Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8]
  wire  _T_1115 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.RocketConfig.fir 294186:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 294188:8 Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 294188:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 294188:8 Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 294188:8]
  wire  _T_1117 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.RocketConfig.fir 294188:8]
  wire  _T_1118 = _T_1115 | _T_1117; // @[Monitor.scala 689:72 chipyard.TestHarness.RocketConfig.fir 294189:8]
  wire  _T_1120 = _T_1118 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294191:8]
  wire  _T_1121 = ~_T_1120; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294192:8]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.RocketConfig.fir 294037:4 Monitor.scala 638:19 chipyard.TestHarness.RocketConfig.fir 294047:4]
  wire [7:0] _GEN_80 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.RocketConfig.fir 294197:8]
  wire  _T_1122 = _GEN_80 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.RocketConfig.fir 294197:8]
  wire  _T_1124 = _T_1122 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294199:8]
  wire  _T_1125 = ~_T_1124; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294200:8]
  wire  _T_1127 = _T_1085 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.RocketConfig.fir 294208:4]
  wire  _T_1128 = _T_1127 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.RocketConfig.fir 294209:4]
  wire  _T_1130 = _T_1128 & _source_ok_T_1; // @[Monitor.scala 694:65 chipyard.TestHarness.RocketConfig.fir 294211:4]
  wire  _T_1132 = _T_1130 & _T_1087; // @[Monitor.scala 694:116 chipyard.TestHarness.RocketConfig.fir 294213:4]
  wire  _T_1133 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.RocketConfig.fir 294215:6]
  wire  _T_1134 = _T_1133 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.RocketConfig.fir 294216:6]
  wire  _T_1136 = _T_1134 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294218:6]
  wire  _T_1137 = ~_T_1136; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294219:6]
  wire  a_set_wo_ready = _GEN_15[0]; // @[chipyard.TestHarness.RocketConfig.fir 294020:4]
  wire  d_clr_wo_ready = _GEN_21[0]; // @[chipyard.TestHarness.RocketConfig.fir 294107:4]
  wire  _T_1138 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.RocketConfig.fir 294225:4]
  wire  _T_1139 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.RocketConfig.fir 294226:4]
  wire  _T_1140 = ~_T_1139; // @[Monitor.scala 699:51 chipyard.TestHarness.RocketConfig.fir 294227:4]
  wire  _T_1141 = _T_1138 | _T_1140; // @[Monitor.scala 699:48 chipyard.TestHarness.RocketConfig.fir 294228:4]
  wire  _T_1143 = _T_1141 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294230:4]
  wire  _T_1144 = ~_T_1143; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294231:4]
  wire  a_set = _GEN_16[0]; // @[chipyard.TestHarness.RocketConfig.fir 294018:4]
  wire  _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.RocketConfig.fir 294236:4]
  wire  d_clr = _GEN_22[0]; // @[chipyard.TestHarness.RocketConfig.fir 294105:4]
  wire  _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.RocketConfig.fir 294237:4]
  wire  _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.RocketConfig.fir 294238:4]
  wire [3:0] a_opcodes_set = _GEN_19[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 294022:4]
  wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.RocketConfig.fir 294240:4]
  wire [3:0] d_opcodes_clr = _GEN_23[3:0]; // @[chipyard.TestHarness.RocketConfig.fir 294109:4]
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.RocketConfig.fir 294241:4]
  wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.RocketConfig.fir 294242:4]
  wire [7:0] a_sizes_set = _GEN_20[7:0]; // @[chipyard.TestHarness.RocketConfig.fir 294024:4]
  wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.RocketConfig.fir 294244:4]
  wire [7:0] d_sizes_clr = _GEN_24[7:0]; // @[chipyard.TestHarness.RocketConfig.fir 294111:4]
  wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56 chipyard.TestHarness.RocketConfig.fir 294245:4]
  wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.RocketConfig.fir 294246:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 294248:4]
  wire  _T_1145 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.RocketConfig.fir 294251:4]
  wire  _T_1146 = ~_T_1145; // @[Monitor.scala 709:16 chipyard.TestHarness.RocketConfig.fir 294252:4]
  wire  _T_1147 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.RocketConfig.fir 294253:4]
  wire  _T_1148 = _T_1146 | _T_1147; // @[Monitor.scala 709:30 chipyard.TestHarness.RocketConfig.fir 294254:4]
  wire  _T_1149 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.RocketConfig.fir 294255:4]
  wire  _T_1150 = _T_1148 | _T_1149; // @[Monitor.scala 709:47 chipyard.TestHarness.RocketConfig.fir 294256:4]
  wire  _T_1152 = _T_1150 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 294258:4]
  wire  _T_1153 = ~_T_1152; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 294259:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.RocketConfig.fir 294265:4]
  wire  _T_1156 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.RocketConfig.fir 294269:4]
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 294275:4]
  reg [8:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 294310:4]
  wire [8:0] d_first_counter1_2 = d_first_counter_2 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.RocketConfig.fir 294312:4]
  wire  d_first_2 = d_first_counter_2 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.RocketConfig.fir 294313:4]
  wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.RocketConfig.fir 294346:4]
  wire [15:0] _GEN_84 = {{8'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.RocketConfig.fir 294351:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_84 & _a_size_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.RocketConfig.fir 294351:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.RocketConfig.fir 294352:4]
  wire  _T_1174 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.RocketConfig.fir 294430:4]
  wire  _T_1176 = _T_1174 & _T_881; // @[Monitor.scala 779:71 chipyard.TestHarness.RocketConfig.fir 294432:4]
  wire  _T_1178 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.RocketConfig.fir 294438:4]
  wire  _T_1180 = _T_1178 & _T_881; // @[Monitor.scala 783:72 chipyard.TestHarness.RocketConfig.fir 294440:4]
  wire [30:0] _GEN_69 = _T_1180 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.RocketConfig.fir 294441:4 Monitor.scala 786:21 chipyard.TestHarness.RocketConfig.fir 294457:6 chipyard.TestHarness.RocketConfig.fir 294428:4]
  wire  _T_1184 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.RocketConfig.fir 294476:6]
  wire  _T_1188 = _T_1184 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294480:6]
  wire  _T_1189 = ~_T_1188; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294481:6]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.RocketConfig.fir 294334:4 Monitor.scala 747:21 chipyard.TestHarness.RocketConfig.fir 294353:4]
  wire  _T_1194 = _GEN_80 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.RocketConfig.fir 294499:8]
  wire  _T_1196 = _T_1194 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294501:8]
  wire  _T_1197 = ~_T_1196; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294502:8]
  wire [7:0] d_sizes_clr_1 = _GEN_69[7:0]; // @[chipyard.TestHarness.RocketConfig.fir 294427:4]
  wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58 chipyard.TestHarness.RocketConfig.fir 294552:4]
  wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.RocketConfig.fir 294553:4]
  wire  _GEN_90 = io_in_a_valid & _T_15; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292482:10]
  wire  _GEN_100 = io_in_a_valid & _T_171; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292672:10]
  wire  _GEN_112 = io_in_a_valid & _T_331; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292810:10]
  wire  _GEN_120 = io_in_a_valid & _T_426; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293002:10]
  wire  _GEN_126 = io_in_a_valid & _T_517; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293115:10]
  wire  _GEN_132 = io_in_a_valid & _T_610; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293225:10]
  wire  _GEN_138 = io_in_a_valid & _T_696; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293333:10]
  wire  _GEN_144 = io_in_a_valid & _T_782; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293446:10]
  wire  _GEN_150 = io_in_d_valid & _T_881; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293509:10]
  wire  _GEN_160 = io_in_d_valid & _T_901; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293551:10]
  wire  _GEN_170 = io_in_d_valid & _T_929; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293609:10]
  wire  _GEN_180 = io_in_d_valid & _T_958; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293668:10]
  wire  _GEN_186 = io_in_d_valid & _T_975; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293703:10]
  wire  _GEN_192 = io_in_d_valid & _T_993; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293739:10]
  wire  _GEN_198 = _T_1088 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294172:10]
  wire  _GEN_203 = _T_1088 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294194:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 294249:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 294556:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 293808:4]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 293808:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 293818:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 293819:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 293807:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 293873:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.RocketConfig.fir 293874:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 293873:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.RocketConfig.fir 293876:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.RocketConfig.fir 293873:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.RocketConfig.fir 293878:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 293888:4]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 293888:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 293898:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 293899:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 293887:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 293962:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.RocketConfig.fir 293963:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 293962:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.RocketConfig.fir 293964:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 293962:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.RocketConfig.fir 293965:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 293962:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.RocketConfig.fir 293966:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 293962:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.RocketConfig.fir 293967:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.RocketConfig.fir 293962:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.RocketConfig.fir 293968:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 293970:4]
      inflight <= 1'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.RocketConfig.fir 293970:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.RocketConfig.fir 294239:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 293971:4]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.RocketConfig.fir 293971:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.RocketConfig.fir 294243:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 293972:4]
      inflight_sizes <= 8'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.RocketConfig.fir 293972:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.RocketConfig.fir 294247:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 293982:4]
      a_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 293982:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 293992:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 293993:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 293807:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 9'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 294004:4]
      d_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 294004:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 294014:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 294015:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 293887:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 9'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 294248:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.RocketConfig.fir 294248:4]
    end else if (_T_1156) begin // @[Monitor.scala 712:47 chipyard.TestHarness.RocketConfig.fir 294270:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.RocketConfig.fir 294271:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.RocketConfig.fir 294266:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 294275:4]
      inflight_sizes_1 <= 8'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.RocketConfig.fir 294275:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.RocketConfig.fir 294554:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 294310:4]
      d_first_counter_2 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.RocketConfig.fir 294310:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.RocketConfig.fir 294320:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.RocketConfig.fir 294321:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.RocketConfig.fir 293887:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 9'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_15 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292482:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292483:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292549:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292550:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292564:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292565:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292571:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292572:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292588:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292589:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292672:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292673:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292739:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292740:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292754:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292755:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292761:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292762:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292777:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292778:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292786:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292787:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_331 & _T_340) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292810:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_340) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292811:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_407) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292881:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_407) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292882:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292895:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292896:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292911:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 292912:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_426 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293002:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293003:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_120 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293016:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293017:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_120 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293032:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293033:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_517 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293115:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293116:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_126 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293129:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293130:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_126 & _T_609) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293147:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_609) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293148:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_610 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293225:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293226:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293239:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293240:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293255:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293256:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_696 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293333:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293334:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293347:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293348:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293363:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293364:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_782 & _T_858) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293446:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_858) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293447:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293460:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293461:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293476:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293477:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293495:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293496:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_881 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293509:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293510:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293517:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293518:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293525:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293526:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293533:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293534:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_900) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293541:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_900) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293542:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_901 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293551:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293552:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293566:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293567:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293574:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293575:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293582:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293583:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293590:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293591:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_929 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293609:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293610:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293624:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293625:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293632:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293633:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293640:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293641:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293649:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293650:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_958 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293668:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293669:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_180 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293676:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293677:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_180 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293684:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293685:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_975 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293703:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293704:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293711:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293712:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293720:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293721:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_993 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293739:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293740:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_192 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293747:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293748:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_192 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293755:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293756:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293835:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293836:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293851:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293852:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293867:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 293868:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293916:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293917:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293924:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293925:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293932:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293933:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293940:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293941:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293948:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293949:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293956:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 293957:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 294101:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 294102:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294161:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294162:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & same_cycle_resp & _T_1109) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294172:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_1109) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294173:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_1113) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294180:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_1113) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294181:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & ~same_cycle_resp & _T_1121) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294194:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_1121) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294195:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_1125) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294202:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_1125) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294203:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294221:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294222:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1144) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 8 (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294233:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1144) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294234:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1153) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 294261:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1153) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.RocketConfig.fir 294262:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294483:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294484:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294504:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.RocketConfig.fir 294505:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  address = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  d_first_counter = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  opcode_1 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  param_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  size_1 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  source_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sink = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  denied = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inflight = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inflight_opcodes = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  inflight_sizes = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_14[8:0];
  _RAND_15 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  watchdog = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_21_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 294711:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 294712:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 294713:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input  [3:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input  [31:0] auto_in_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output [3:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output        auto_out_a_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output [31:0] auto_out_a_bits_address, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input  [3:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input         auto_out_d_bits_source, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input  [2:0]  auto_out_d_bits_sink, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.RocketConfig.fir 294714:4]
);
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire [2:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [31:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire  bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [31:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire  bundleOut_0_a_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire [1:0] bundleIn_0_d_q_io_enq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire [3:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_io_enq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_io_enq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire [3:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
  TLMonitor_57_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.RocketConfig.fir 294721:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_6_inTestHarness bundleOut_0_a_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294748:4]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
  );
  Queue_7_inTestHarness bundleIn_0_d_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.RocketConfig.fir 294762:4]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
    .io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Decoupled.scala 299:17 chipyard.TestHarness.RocketConfig.fir 294760:4]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 294775:4]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 294775:4]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 294761:4]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 294761:4]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 294761:4]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 294761:4]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 294761:4]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 294761:4]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 294761:4]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 294761:4]
  assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 Buffer.scala 37:13 chipyard.TestHarness.RocketConfig.fir 294761:4]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 Decoupled.scala 299:17 chipyard.TestHarness.RocketConfig.fir 294774:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 294722:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 294723:4]
  assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Decoupled.scala 299:17 chipyard.TestHarness.RocketConfig.fir 294760:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 294775:4]
  assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 294775:4]
  assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 294775:4]
  assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 294775:4]
  assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 294775:4]
  assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 294775:4]
  assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 294775:4]
  assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 Buffer.scala 38:13 chipyard.TestHarness.RocketConfig.fir 294775:4]
  assign bundleOut_0_a_q_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 294749:4]
  assign bundleOut_0_a_q_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 294750:4]
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 294746:4]
  assign bundleIn_0_d_q_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 294763:4]
  assign bundleIn_0_d_q_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 294764:4]
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 294746:4]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 294746:4]
  assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 294746:4]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 294746:4]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 294746:4]
  assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 294746:4]
  assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 294746:4]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 294746:4]
  assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.RocketConfig.fir 294744:4 LazyModule.scala 311:12 chipyard.TestHarness.RocketConfig.fir 294746:4]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.RocketConfig.fir 294719:4 LazyModule.scala 309:16 chipyard.TestHarness.RocketConfig.fir 294747:4]
endmodule
module SerialRAM_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 294795:2]
  input         clock, // @[chipyard.TestHarness.RocketConfig.fir 294796:4]
  input         reset, // @[chipyard.TestHarness.RocketConfig.fir 294797:4]
  input         io_ser_in_ready, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  output        io_ser_in_valid, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  output [3:0]  io_ser_in_bits, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  output        io_ser_out_ready, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  input         io_ser_out_valid, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  input  [3:0]  io_ser_out_bits, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  output        io_tsi_ser_in_ready, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  input         io_tsi_ser_in_valid, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  input  [31:0] io_tsi_ser_in_bits, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  input         io_tsi_ser_out_ready, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  output        io_tsi_ser_out_valid, // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
  output [31:0] io_tsi_ser_out_bits // @[chipyard.TestHarness.RocketConfig.fir 294799:4]
);
  wire  adapter_clock; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire  adapter_reset; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire  adapter_auto_out_a_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire  adapter_auto_out_a_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire [2:0] adapter_auto_out_a_bits_opcode; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire [3:0] adapter_auto_out_a_bits_size; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire [31:0] adapter_auto_out_a_bits_address; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire [7:0] adapter_auto_out_a_bits_mask; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire [63:0] adapter_auto_out_a_bits_data; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire  adapter_auto_out_d_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire  adapter_auto_out_d_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire [63:0] adapter_auto_out_d_bits_data; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire  adapter_io_serial_in_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire  adapter_io_serial_in_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire [31:0] adapter_io_serial_in_bits; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire  adapter_io_serial_out_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire  adapter_io_serial_out_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire [31:0] adapter_io_serial_out_bits; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
  wire  serdesser_clock; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_reset; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_manager_in_a_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_manager_in_a_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [2:0] serdesser_auto_manager_in_a_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [2:0] serdesser_auto_manager_in_a_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [3:0] serdesser_auto_manager_in_a_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_manager_in_a_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [31:0] serdesser_auto_manager_in_a_bits_address; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [7:0] serdesser_auto_manager_in_a_bits_mask; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [63:0] serdesser_auto_manager_in_a_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_manager_in_a_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_manager_in_d_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_manager_in_d_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [2:0] serdesser_auto_manager_in_d_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [1:0] serdesser_auto_manager_in_d_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [3:0] serdesser_auto_manager_in_d_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_manager_in_d_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [2:0] serdesser_auto_manager_in_d_bits_sink; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_manager_in_d_bits_denied; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [63:0] serdesser_auto_manager_in_d_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_manager_in_d_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_client_out_a_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_client_out_a_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [2:0] serdesser_auto_client_out_a_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [2:0] serdesser_auto_client_out_a_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [2:0] serdesser_auto_client_out_a_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [3:0] serdesser_auto_client_out_a_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [28:0] serdesser_auto_client_out_a_bits_address; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [7:0] serdesser_auto_client_out_a_bits_mask; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [63:0] serdesser_auto_client_out_a_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_client_out_a_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_client_out_d_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_client_out_d_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [2:0] serdesser_auto_client_out_d_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [1:0] serdesser_auto_client_out_d_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [2:0] serdesser_auto_client_out_d_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [3:0] serdesser_auto_client_out_d_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_client_out_d_bits_sink; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_client_out_d_bits_denied; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [63:0] serdesser_auto_client_out_d_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_auto_client_out_d_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_io_ser_in_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_io_ser_in_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [3:0] serdesser_io_ser_in_bits; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_io_ser_out_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  serdesser_io_ser_out_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire [3:0] serdesser_io_ser_out_bits; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
  wire  srams_clock; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire  srams_reset; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire  srams_auto_in_a_ready; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire  srams_auto_in_a_valid; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [2:0] srams_auto_in_a_bits_opcode; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [2:0] srams_auto_in_a_bits_param; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [1:0] srams_auto_in_a_bits_size; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [7:0] srams_auto_in_a_bits_source; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [28:0] srams_auto_in_a_bits_address; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [7:0] srams_auto_in_a_bits_mask; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [63:0] srams_auto_in_a_bits_data; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire  srams_auto_in_a_bits_corrupt; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire  srams_auto_in_d_ready; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire  srams_auto_in_d_valid; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [2:0] srams_auto_in_d_bits_opcode; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [1:0] srams_auto_in_d_bits_size; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [7:0] srams_auto_in_d_bits_source; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire [63:0] srams_auto_in_d_bits_data; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
  wire  xbar_auto_in_a_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_in_a_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [2:0] xbar_auto_in_a_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [2:0] xbar_auto_in_a_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [2:0] xbar_auto_in_a_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [3:0] xbar_auto_in_a_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [28:0] xbar_auto_in_a_bits_address; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [7:0] xbar_auto_in_a_bits_mask; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [63:0] xbar_auto_in_a_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_in_a_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_in_d_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_in_d_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [2:0] xbar_auto_in_d_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [1:0] xbar_auto_in_d_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [2:0] xbar_auto_in_d_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [3:0] xbar_auto_in_d_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_in_d_bits_sink; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_in_d_bits_denied; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [63:0] xbar_auto_in_d_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_in_d_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_out_a_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_out_a_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [2:0] xbar_auto_out_a_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [2:0] xbar_auto_out_a_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [2:0] xbar_auto_out_a_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [3:0] xbar_auto_out_a_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [28:0] xbar_auto_out_a_bits_address; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [7:0] xbar_auto_out_a_bits_mask; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [63:0] xbar_auto_out_a_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_out_a_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_out_d_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_out_d_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [2:0] xbar_auto_out_d_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [1:0] xbar_auto_out_d_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [2:0] xbar_auto_out_d_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [3:0] xbar_auto_out_d_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_out_d_bits_sink; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_out_d_bits_denied; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire [63:0] xbar_auto_out_d_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  xbar_auto_out_d_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
  wire  buffer_clock; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_reset; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [1:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [7:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [28:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_in_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [1:0] buffer_auto_in_d_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [1:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [7:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_in_d_bits_sink; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [1:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [7:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [28:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_out_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [1:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [7:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [2:0] fragmenter_auto_in_a_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [2:0] fragmenter_auto_in_a_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [3:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [28:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [7:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [63:0] fragmenter_auto_in_a_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_in_a_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [2:0] fragmenter_auto_in_d_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [1:0] fragmenter_auto_in_d_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [3:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_in_d_bits_sink; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_in_d_bits_denied; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [63:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_in_d_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [2:0] fragmenter_auto_out_a_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [2:0] fragmenter_auto_out_a_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [7:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [28:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [7:0] fragmenter_auto_out_a_bits_mask; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [63:0] fragmenter_auto_out_a_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_out_a_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [2:0] fragmenter_auto_out_d_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [1:0] fragmenter_auto_out_d_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [7:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_out_d_bits_sink; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_out_d_bits_denied; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire [63:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  fragmenter_auto_out_d_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
  wire  buffer_1_clock; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_reset; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_in_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_in_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [2:0] buffer_1_auto_in_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [3:0] buffer_1_auto_in_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [31:0] buffer_1_auto_in_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [7:0] buffer_1_auto_in_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [63:0] buffer_1_auto_in_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_in_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_in_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [63:0] buffer_1_auto_in_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_out_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_out_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [2:0] buffer_1_auto_out_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [2:0] buffer_1_auto_out_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [3:0] buffer_1_auto_out_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_out_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [31:0] buffer_1_auto_out_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [7:0] buffer_1_auto_out_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [63:0] buffer_1_auto_out_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_out_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_out_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_out_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [2:0] buffer_1_auto_out_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [1:0] buffer_1_auto_out_d_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [3:0] buffer_1_auto_out_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_out_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [2:0] buffer_1_auto_out_d_bits_sink; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_out_d_bits_denied; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire [63:0] buffer_1_auto_out_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  wire  buffer_1_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
  SerialAdapter_inTestHarness adapter ( // @[SerialAdapter.scala 311:27 chipyard.TestHarness.RocketConfig.fir 294805:4]
    .clock(adapter_clock),
    .reset(adapter_reset),
    .auto_out_a_ready(adapter_auto_out_a_ready),
    .auto_out_a_valid(adapter_auto_out_a_valid),
    .auto_out_a_bits_opcode(adapter_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(adapter_auto_out_a_bits_size),
    .auto_out_a_bits_address(adapter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(adapter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(adapter_auto_out_a_bits_data),
    .auto_out_d_ready(adapter_auto_out_d_ready),
    .auto_out_d_valid(adapter_auto_out_d_valid),
    .auto_out_d_bits_data(adapter_auto_out_d_bits_data),
    .io_serial_in_ready(adapter_io_serial_in_ready),
    .io_serial_in_valid(adapter_io_serial_in_valid),
    .io_serial_in_bits(adapter_io_serial_in_bits),
    .io_serial_out_ready(adapter_io_serial_out_ready),
    .io_serial_out_valid(adapter_io_serial_out_valid),
    .io_serial_out_bits(adapter_io_serial_out_bits)
  );
  TLSerdesser_1_inTestHarness serdesser ( // @[SerialAdapter.scala 312:29 chipyard.TestHarness.RocketConfig.fir 294812:4]
    .clock(serdesser_clock),
    .reset(serdesser_reset),
    .auto_manager_in_a_ready(serdesser_auto_manager_in_a_ready),
    .auto_manager_in_a_valid(serdesser_auto_manager_in_a_valid),
    .auto_manager_in_a_bits_opcode(serdesser_auto_manager_in_a_bits_opcode),
    .auto_manager_in_a_bits_param(serdesser_auto_manager_in_a_bits_param),
    .auto_manager_in_a_bits_size(serdesser_auto_manager_in_a_bits_size),
    .auto_manager_in_a_bits_source(serdesser_auto_manager_in_a_bits_source),
    .auto_manager_in_a_bits_address(serdesser_auto_manager_in_a_bits_address),
    .auto_manager_in_a_bits_mask(serdesser_auto_manager_in_a_bits_mask),
    .auto_manager_in_a_bits_data(serdesser_auto_manager_in_a_bits_data),
    .auto_manager_in_a_bits_corrupt(serdesser_auto_manager_in_a_bits_corrupt),
    .auto_manager_in_d_ready(serdesser_auto_manager_in_d_ready),
    .auto_manager_in_d_valid(serdesser_auto_manager_in_d_valid),
    .auto_manager_in_d_bits_opcode(serdesser_auto_manager_in_d_bits_opcode),
    .auto_manager_in_d_bits_param(serdesser_auto_manager_in_d_bits_param),
    .auto_manager_in_d_bits_size(serdesser_auto_manager_in_d_bits_size),
    .auto_manager_in_d_bits_source(serdesser_auto_manager_in_d_bits_source),
    .auto_manager_in_d_bits_sink(serdesser_auto_manager_in_d_bits_sink),
    .auto_manager_in_d_bits_denied(serdesser_auto_manager_in_d_bits_denied),
    .auto_manager_in_d_bits_data(serdesser_auto_manager_in_d_bits_data),
    .auto_manager_in_d_bits_corrupt(serdesser_auto_manager_in_d_bits_corrupt),
    .auto_client_out_a_ready(serdesser_auto_client_out_a_ready),
    .auto_client_out_a_valid(serdesser_auto_client_out_a_valid),
    .auto_client_out_a_bits_opcode(serdesser_auto_client_out_a_bits_opcode),
    .auto_client_out_a_bits_param(serdesser_auto_client_out_a_bits_param),
    .auto_client_out_a_bits_size(serdesser_auto_client_out_a_bits_size),
    .auto_client_out_a_bits_source(serdesser_auto_client_out_a_bits_source),
    .auto_client_out_a_bits_address(serdesser_auto_client_out_a_bits_address),
    .auto_client_out_a_bits_mask(serdesser_auto_client_out_a_bits_mask),
    .auto_client_out_a_bits_data(serdesser_auto_client_out_a_bits_data),
    .auto_client_out_a_bits_corrupt(serdesser_auto_client_out_a_bits_corrupt),
    .auto_client_out_d_ready(serdesser_auto_client_out_d_ready),
    .auto_client_out_d_valid(serdesser_auto_client_out_d_valid),
    .auto_client_out_d_bits_opcode(serdesser_auto_client_out_d_bits_opcode),
    .auto_client_out_d_bits_param(serdesser_auto_client_out_d_bits_param),
    .auto_client_out_d_bits_size(serdesser_auto_client_out_d_bits_size),
    .auto_client_out_d_bits_source(serdesser_auto_client_out_d_bits_source),
    .auto_client_out_d_bits_sink(serdesser_auto_client_out_d_bits_sink),
    .auto_client_out_d_bits_denied(serdesser_auto_client_out_d_bits_denied),
    .auto_client_out_d_bits_data(serdesser_auto_client_out_d_bits_data),
    .auto_client_out_d_bits_corrupt(serdesser_auto_client_out_d_bits_corrupt),
    .io_ser_in_ready(serdesser_io_ser_in_ready),
    .io_ser_in_valid(serdesser_io_ser_in_valid),
    .io_ser_in_bits(serdesser_io_ser_in_bits),
    .io_ser_out_ready(serdesser_io_ser_out_ready),
    .io_ser_out_valid(serdesser_io_ser_out_valid),
    .io_ser_out_bits(serdesser_io_ser_out_bits)
  );
  TLRAM_inTestHarness srams ( // @[SerialAdapter.scala 322:15 chipyard.TestHarness.RocketConfig.fir 294819:4]
    .clock(srams_clock),
    .reset(srams_reset),
    .auto_in_a_ready(srams_auto_in_a_ready),
    .auto_in_a_valid(srams_auto_in_a_valid),
    .auto_in_a_bits_opcode(srams_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(srams_auto_in_a_bits_param),
    .auto_in_a_bits_size(srams_auto_in_a_bits_size),
    .auto_in_a_bits_source(srams_auto_in_a_bits_source),
    .auto_in_a_bits_address(srams_auto_in_a_bits_address),
    .auto_in_a_bits_mask(srams_auto_in_a_bits_mask),
    .auto_in_a_bits_data(srams_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(srams_auto_in_a_bits_corrupt),
    .auto_in_d_ready(srams_auto_in_d_ready),
    .auto_in_d_valid(srams_auto_in_d_valid),
    .auto_in_d_bits_opcode(srams_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(srams_auto_in_d_bits_size),
    .auto_in_d_bits_source(srams_auto_in_d_bits_source),
    .auto_in_d_bits_data(srams_auto_in_d_bits_data)
  );
  TLXbar_10_inTestHarness xbar ( // @[Xbar.scala 142:26 chipyard.TestHarness.RocketConfig.fir 294825:4]
    .auto_in_a_ready(xbar_auto_in_a_ready),
    .auto_in_a_valid(xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(xbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(xbar_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(xbar_auto_in_a_bits_corrupt),
    .auto_in_d_ready(xbar_auto_in_d_ready),
    .auto_in_d_valid(xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(xbar_auto_in_d_bits_param),
    .auto_in_d_bits_size(xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(xbar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(xbar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(xbar_auto_in_d_bits_corrupt),
    .auto_out_a_ready(xbar_auto_out_a_ready),
    .auto_out_a_valid(xbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(xbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(xbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(xbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(xbar_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(xbar_auto_out_a_bits_corrupt),
    .auto_out_d_ready(xbar_auto_out_d_ready),
    .auto_out_d_valid(xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(xbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(xbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(xbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(xbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(xbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(xbar_auto_out_d_bits_corrupt)
  );
  TLBuffer_20_inTestHarness buffer ( // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294831:4]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data)
  );
  TLFragmenter_8_inTestHarness fragmenter ( // @[Fragmenter.scala 333:34 chipyard.TestHarness.RocketConfig.fir 294837:4]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(fragmenter_auto_in_d_bits_param),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_sink(fragmenter_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(fragmenter_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fragmenter_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(fragmenter_auto_out_d_bits_param),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_sink(fragmenter_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(fragmenter_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fragmenter_auto_out_d_bits_corrupt)
  );
  TLBuffer_21_inTestHarness buffer_1 ( // @[Buffer.scala 68:28 chipyard.TestHarness.RocketConfig.fir 294843:4]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_a_ready(buffer_1_auto_in_a_ready),
    .auto_in_a_valid(buffer_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
    .auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_1_auto_in_d_ready),
    .auto_in_d_valid(buffer_1_auto_in_d_valid),
    .auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
    .auto_out_a_ready(buffer_1_auto_out_a_ready),
    .auto_out_a_valid(buffer_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_1_auto_out_a_bits_corrupt),
    .auto_out_d_ready(buffer_1_auto_out_d_ready),
    .auto_out_d_valid(buffer_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
  );
  assign io_ser_in_valid = serdesser_io_ser_out_valid; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.RocketConfig.fir 294859:4]
  assign io_ser_in_bits = serdesser_io_ser_out_bits; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.RocketConfig.fir 294858:4]
  assign io_ser_out_ready = serdesser_io_ser_in_ready; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.RocketConfig.fir 294857:4]
  assign io_tsi_ser_in_ready = adapter_io_serial_in_ready; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.RocketConfig.fir 294866:4]
  assign io_tsi_ser_out_valid = adapter_io_serial_out_valid; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.RocketConfig.fir 294862:4]
  assign io_tsi_ser_out_bits = adapter_io_serial_out_bits; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.RocketConfig.fir 294861:4]
  assign adapter_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 294810:4]
  assign adapter_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 294811:4]
  assign adapter_auto_out_a_ready = buffer_1_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294849:4]
  assign adapter_auto_out_d_valid = buffer_1_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294849:4]
  assign adapter_auto_out_d_bits_data = buffer_1_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294849:4]
  assign adapter_io_serial_in_valid = io_tsi_ser_in_valid; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.RocketConfig.fir 294865:4]
  assign adapter_io_serial_in_bits = io_tsi_ser_in_bits; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.RocketConfig.fir 294864:4]
  assign adapter_io_serial_out_ready = io_tsi_ser_out_ready; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.RocketConfig.fir 294863:4]
  assign serdesser_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 294817:4]
  assign serdesser_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 294818:4]
  assign serdesser_auto_manager_in_a_valid = buffer_1_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign serdesser_auto_manager_in_a_bits_opcode = buffer_1_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign serdesser_auto_manager_in_a_bits_param = buffer_1_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign serdesser_auto_manager_in_a_bits_size = buffer_1_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign serdesser_auto_manager_in_a_bits_source = buffer_1_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign serdesser_auto_manager_in_a_bits_address = buffer_1_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign serdesser_auto_manager_in_a_bits_mask = buffer_1_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign serdesser_auto_manager_in_a_bits_data = buffer_1_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign serdesser_auto_manager_in_a_bits_corrupt = buffer_1_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign serdesser_auto_manager_in_d_ready = buffer_1_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign serdesser_auto_client_out_a_ready = xbar_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign serdesser_auto_client_out_d_valid = xbar_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign serdesser_auto_client_out_d_bits_opcode = xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign serdesser_auto_client_out_d_bits_param = xbar_auto_in_d_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign serdesser_auto_client_out_d_bits_size = xbar_auto_in_d_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign serdesser_auto_client_out_d_bits_source = xbar_auto_in_d_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign serdesser_auto_client_out_d_bits_sink = xbar_auto_in_d_bits_sink; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign serdesser_auto_client_out_d_bits_denied = xbar_auto_in_d_bits_denied; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign serdesser_auto_client_out_d_bits_data = xbar_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign serdesser_auto_client_out_d_bits_corrupt = xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign serdesser_io_ser_in_valid = io_ser_out_valid; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.RocketConfig.fir 294856:4]
  assign serdesser_io_ser_in_bits = io_ser_out_bits; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.RocketConfig.fir 294855:4]
  assign serdesser_io_ser_out_ready = io_ser_in_ready; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.RocketConfig.fir 294860:4]
  assign srams_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 294823:4]
  assign srams_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 294824:4]
  assign srams_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign srams_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign srams_auto_in_a_bits_param = buffer_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign srams_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign srams_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign srams_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign srams_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign srams_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign srams_auto_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign srams_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign xbar_auto_in_a_valid = serdesser_auto_client_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign xbar_auto_in_a_bits_opcode = serdesser_auto_client_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign xbar_auto_in_a_bits_param = serdesser_auto_client_out_a_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign xbar_auto_in_a_bits_size = serdesser_auto_client_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign xbar_auto_in_a_bits_source = serdesser_auto_client_out_a_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign xbar_auto_in_a_bits_address = serdesser_auto_client_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign xbar_auto_in_a_bits_mask = serdesser_auto_client_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign xbar_auto_in_a_bits_data = serdesser_auto_client_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign xbar_auto_in_a_bits_corrupt = serdesser_auto_client_out_a_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign xbar_auto_in_d_ready = serdesser_auto_client_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294850:4]
  assign xbar_auto_out_a_ready = fragmenter_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign xbar_auto_out_d_valid = fragmenter_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign xbar_auto_out_d_bits_opcode = fragmenter_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign xbar_auto_out_d_bits_param = fragmenter_auto_in_d_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign xbar_auto_out_d_bits_size = fragmenter_auto_in_d_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign xbar_auto_out_d_bits_source = fragmenter_auto_in_d_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign xbar_auto_out_d_bits_sink = fragmenter_auto_in_d_bits_sink; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign xbar_auto_out_d_bits_denied = fragmenter_auto_in_d_bits_denied; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign xbar_auto_out_d_bits_data = fragmenter_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign xbar_auto_out_d_bits_corrupt = fragmenter_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign buffer_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 294835:4]
  assign buffer_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 294836:4]
  assign buffer_auto_in_a_valid = fragmenter_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_auto_in_a_bits_opcode = fragmenter_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_auto_in_a_bits_param = fragmenter_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_auto_in_a_bits_size = fragmenter_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_auto_in_a_bits_source = fragmenter_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_auto_in_a_bits_address = fragmenter_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_auto_in_a_bits_mask = fragmenter_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_auto_in_a_bits_data = fragmenter_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_auto_in_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_auto_in_d_ready = fragmenter_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_auto_out_a_ready = srams_auto_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign buffer_auto_out_d_valid = srams_auto_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign buffer_auto_out_d_bits_opcode = srams_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign buffer_auto_out_d_bits_size = srams_auto_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign buffer_auto_out_d_bits_source = srams_auto_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign buffer_auto_out_d_bits_data = srams_auto_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294852:4]
  assign fragmenter_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 294841:4]
  assign fragmenter_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 294842:4]
  assign fragmenter_auto_in_a_valid = xbar_auto_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign fragmenter_auto_in_a_bits_opcode = xbar_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign fragmenter_auto_in_a_bits_param = xbar_auto_out_a_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign fragmenter_auto_in_a_bits_size = xbar_auto_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign fragmenter_auto_in_a_bits_source = xbar_auto_out_a_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign fragmenter_auto_in_a_bits_address = xbar_auto_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign fragmenter_auto_in_a_bits_mask = xbar_auto_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign fragmenter_auto_in_a_bits_data = xbar_auto_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign fragmenter_auto_in_a_bits_corrupt = xbar_auto_out_a_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign fragmenter_auto_in_d_ready = xbar_auto_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294851:4]
  assign fragmenter_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign fragmenter_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign fragmenter_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign fragmenter_auto_out_d_bits_param = buffer_auto_in_d_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign fragmenter_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign fragmenter_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign fragmenter_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign fragmenter_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign fragmenter_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign fragmenter_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294853:4]
  assign buffer_1_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 294847:4]
  assign buffer_1_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 294848:4]
  assign buffer_1_auto_in_a_valid = adapter_auto_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294849:4]
  assign buffer_1_auto_in_a_bits_opcode = adapter_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294849:4]
  assign buffer_1_auto_in_a_bits_size = adapter_auto_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294849:4]
  assign buffer_1_auto_in_a_bits_address = adapter_auto_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294849:4]
  assign buffer_1_auto_in_a_bits_mask = adapter_auto_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294849:4]
  assign buffer_1_auto_in_a_bits_data = adapter_auto_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294849:4]
  assign buffer_1_auto_in_d_ready = adapter_auto_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.RocketConfig.fir 294849:4]
  assign buffer_1_auto_out_a_ready = serdesser_auto_manager_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign buffer_1_auto_out_d_valid = serdesser_auto_manager_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign buffer_1_auto_out_d_bits_opcode = serdesser_auto_manager_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign buffer_1_auto_out_d_bits_param = serdesser_auto_manager_in_d_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign buffer_1_auto_out_d_bits_size = serdesser_auto_manager_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign buffer_1_auto_out_d_bits_source = serdesser_auto_manager_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign buffer_1_auto_out_d_bits_sink = serdesser_auto_manager_in_d_bits_sink; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign buffer_1_auto_out_d_bits_denied = serdesser_auto_manager_in_d_bits_denied; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign buffer_1_auto_out_d_bits_data = serdesser_auto_manager_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
  assign buffer_1_auto_out_d_bits_corrupt = serdesser_auto_manager_in_d_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.RocketConfig.fir 294854:4]
endmodule
module Queue_44_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 294889:2]
  input        clock, // @[chipyard.TestHarness.RocketConfig.fir 294890:4]
  input        reset, // @[chipyard.TestHarness.RocketConfig.fir 294891:4]
  output       io_enq_ready, // @[chipyard.TestHarness.RocketConfig.fir 294892:4]
  input        io_enq_valid, // @[chipyard.TestHarness.RocketConfig.fir 294892:4]
  input  [7:0] io_enq_bits, // @[chipyard.TestHarness.RocketConfig.fir 294892:4]
  input        io_deq_ready, // @[chipyard.TestHarness.RocketConfig.fir 294892:4]
  output       io_deq_valid, // @[chipyard.TestHarness.RocketConfig.fir 294892:4]
  output [7:0] io_deq_bits // @[chipyard.TestHarness.RocketConfig.fir 294892:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:127]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 294894:4]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 294894:4]
  wire [6:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 294894:4]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 294894:4]
  wire [6:0] ram_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 294894:4]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 294894:4]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 294894:4]
  reg [6:0] enq_ptr_value; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 294895:4]
  reg [6:0] deq_ptr_value; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 294896:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 294897:4]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33 chipyard.TestHarness.RocketConfig.fir 294898:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.RocketConfig.fir 294899:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.RocketConfig.fir 294900:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.RocketConfig.fir 294901:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 294902:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.RocketConfig.fir 294905:4]
  wire [6:0] _value_T_1 = enq_ptr_value + 7'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 294913:6]
  wire [6:0] _value_T_3 = deq_ptr_value + 7'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 294919:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.RocketConfig.fir 294922:4]
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 294894:4]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.RocketConfig.fir 294928:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.RocketConfig.fir 294926:4]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.RocketConfig.fir 294931:4]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.RocketConfig.fir 294894:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 294895:4]
      enq_ptr_value <= 7'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 294895:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.RocketConfig.fir 294908:4]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 294914:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 294896:4]
      deq_ptr_value <= 7'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 294896:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.RocketConfig.fir 294916:4]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 294920:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 294897:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.RocketConfig.fir 294897:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.RocketConfig.fir 294923:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.RocketConfig.fir 294924:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module UARTAdapter_inTestHarness( // @[chipyard.TestHarness.RocketConfig.fir 294997:2]
  input   clock, // @[chipyard.TestHarness.RocketConfig.fir 294998:4]
  input   reset, // @[chipyard.TestHarness.RocketConfig.fir 294999:4]
  input   io_uart_txd, // @[chipyard.TestHarness.RocketConfig.fir 295000:4]
  output  io_uart_rxd // @[chipyard.TestHarness.RocketConfig.fir 295000:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  txfifo_clock; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.RocketConfig.fir 295002:4]
  wire  txfifo_reset; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.RocketConfig.fir 295002:4]
  wire  txfifo_io_enq_ready; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.RocketConfig.fir 295002:4]
  wire  txfifo_io_enq_valid; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.RocketConfig.fir 295002:4]
  wire [7:0] txfifo_io_enq_bits; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.RocketConfig.fir 295002:4]
  wire  txfifo_io_deq_ready; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.RocketConfig.fir 295002:4]
  wire  txfifo_io_deq_valid; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.RocketConfig.fir 295002:4]
  wire [7:0] txfifo_io_deq_bits; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.RocketConfig.fir 295002:4]
  wire  rxfifo_clock; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.RocketConfig.fir 295005:4]
  wire  rxfifo_reset; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.RocketConfig.fir 295005:4]
  wire  rxfifo_io_enq_ready; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.RocketConfig.fir 295005:4]
  wire  rxfifo_io_enq_valid; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.RocketConfig.fir 295005:4]
  wire [7:0] rxfifo_io_enq_bits; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.RocketConfig.fir 295005:4]
  wire  rxfifo_io_deq_ready; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.RocketConfig.fir 295005:4]
  wire  rxfifo_io_deq_valid; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.RocketConfig.fir 295005:4]
  wire [7:0] rxfifo_io_deq_bits; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.RocketConfig.fir 295005:4]
  wire  sim_clock; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.RocketConfig.fir 295154:4]
  wire  sim_reset; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.RocketConfig.fir 295154:4]
  wire  sim_serial_in_ready; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.RocketConfig.fir 295154:4]
  wire  sim_serial_in_valid; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.RocketConfig.fir 295154:4]
  wire [7:0] sim_serial_in_bits; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.RocketConfig.fir 295154:4]
  wire  sim_serial_out_ready; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.RocketConfig.fir 295154:4]
  wire  sim_serial_out_valid; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.RocketConfig.fir 295154:4]
  wire [7:0] sim_serial_out_bits; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.RocketConfig.fir 295154:4]
  reg [1:0] txState; // @[UARTAdapter.scala 38:24 chipyard.TestHarness.RocketConfig.fir 295008:4]
  reg [7:0] txData; // @[UARTAdapter.scala 39:19 chipyard.TestHarness.RocketConfig.fir 295009:4]
  wire  _T = txState == 2'h2; // @[UARTAdapter.scala 41:49 chipyard.TestHarness.RocketConfig.fir 295010:4]
  wire  _T_1 = _T & txfifo_io_enq_ready; // @[UARTAdapter.scala 41:61 chipyard.TestHarness.RocketConfig.fir 295011:4]
  reg [2:0] txDataIdx; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295012:4]
  wire  wrap_wrap = txDataIdx == 3'h7; // @[Counter.scala 72:24 chipyard.TestHarness.RocketConfig.fir 295016:6]
  wire [2:0] _wrap_value_T_1 = txDataIdx + 3'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 295018:6]
  wire  txDataWrap = _T_1 & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295015:4 Counter.scala 118:24 chipyard.TestHarness.RocketConfig.fir 295020:6 chipyard.TestHarness.RocketConfig.fir 295014:4]
  wire  _T_2 = txState == 2'h1; // @[UARTAdapter.scala 43:51 chipyard.TestHarness.RocketConfig.fir 295022:4]
  wire  _T_3 = _T_2 & txfifo_io_enq_ready; // @[UARTAdapter.scala 43:63 chipyard.TestHarness.RocketConfig.fir 295023:4]
  reg [9:0] txBaudCount; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295024:4]
  wire  wrap_wrap_1 = txBaudCount == 10'h363; // @[Counter.scala 72:24 chipyard.TestHarness.RocketConfig.fir 295028:6]
  wire [9:0] _wrap_value_T_3 = txBaudCount + 10'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 295030:6]
  wire  txBaudWrap = _T_3 & wrap_wrap_1; // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295027:4 Counter.scala 118:24 chipyard.TestHarness.RocketConfig.fir 295035:6 chipyard.TestHarness.RocketConfig.fir 295026:4]
  wire  _T_4 = txState == 2'h0; // @[UARTAdapter.scala 44:53 chipyard.TestHarness.RocketConfig.fir 295037:4]
  wire  _T_5 = ~io_uart_txd; // @[UARTAdapter.scala 44:80 chipyard.TestHarness.RocketConfig.fir 295038:4]
  wire  _T_6 = _T_4 & _T_5; // @[UARTAdapter.scala 44:65 chipyard.TestHarness.RocketConfig.fir 295039:4]
  wire  _T_7 = _T_6 & txfifo_io_enq_ready; // @[UARTAdapter.scala 44:88 chipyard.TestHarness.RocketConfig.fir 295040:4]
  reg [1:0] txSlackCount; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295041:4]
  wire  wrap_wrap_2 = txSlackCount == 2'h3; // @[Counter.scala 72:24 chipyard.TestHarness.RocketConfig.fir 295045:6]
  wire [1:0] _wrap_value_T_5 = txSlackCount + 2'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 295047:6]
  wire  txSlackWrap = _T_7 & wrap_wrap_2; // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295044:4 Counter.scala 118:24 chipyard.TestHarness.RocketConfig.fir 295049:6 chipyard.TestHarness.RocketConfig.fir 295043:4]
  wire  _T_8 = 2'h0 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.RocketConfig.fir 295051:4]
  wire  _T_9 = 2'h1 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.RocketConfig.fir 295059:6]
  wire  _T_10 = 2'h2 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.RocketConfig.fir 295066:8]
  wire [7:0] _GEN_35 = {{7'd0}, io_uart_txd}; // @[UARTAdapter.scala 60:41 chipyard.TestHarness.RocketConfig.fir 295069:12]
  wire [7:0] _txData_T = _GEN_35 << txDataIdx; // @[UARTAdapter.scala 60:41 chipyard.TestHarness.RocketConfig.fir 295069:12]
  wire [7:0] _txData_T_1 = txData | _txData_T; // @[UARTAdapter.scala 60:26 chipyard.TestHarness.RocketConfig.fir 295070:12]
  wire [1:0] _txState_T_1 = io_uart_txd ? 2'h0 : 2'h3; // @[UARTAdapter.scala 63:23 chipyard.TestHarness.RocketConfig.fir 295075:12]
  wire [1:0] _GEN_11 = txfifo_io_enq_ready ? 2'h1 : txState; // @[UARTAdapter.scala 64:39 chipyard.TestHarness.RocketConfig.fir 295079:12 UARTAdapter.scala 65:17 chipyard.TestHarness.RocketConfig.fir 295080:14 UARTAdapter.scala 38:24 chipyard.TestHarness.RocketConfig.fir 295008:4]
  wire [1:0] _GEN_12 = txDataWrap ? _txState_T_1 : _GEN_11; // @[UARTAdapter.scala 62:24 chipyard.TestHarness.RocketConfig.fir 295073:10 UARTAdapter.scala 63:17 chipyard.TestHarness.RocketConfig.fir 295076:12]
  wire  _T_11 = 2'h3 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.RocketConfig.fir 295084:10]
  wire  _T_13 = io_uart_txd & txfifo_io_enq_ready; // @[UARTAdapter.scala 69:32 chipyard.TestHarness.RocketConfig.fir 295087:12]
  wire [1:0] _GEN_13 = _T_13 ? 2'h0 : txState; // @[UARTAdapter.scala 69:56 chipyard.TestHarness.RocketConfig.fir 295088:12 UARTAdapter.scala 70:17 chipyard.TestHarness.RocketConfig.fir 295089:14 UARTAdapter.scala 38:24 chipyard.TestHarness.RocketConfig.fir 295008:4]
  wire [1:0] _GEN_14 = _T_11 ? _GEN_13 : txState; // @[Conditional.scala 39:67 chipyard.TestHarness.RocketConfig.fir 295085:10 UARTAdapter.scala 38:24 chipyard.TestHarness.RocketConfig.fir 295008:4]
  reg [1:0] rxState; // @[UARTAdapter.scala 79:24 chipyard.TestHarness.RocketConfig.fir 295094:4]
  reg [9:0] rxBaudCount; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295095:4]
  wire  wrap_wrap_3 = rxBaudCount == 10'h363; // @[Counter.scala 72:24 chipyard.TestHarness.RocketConfig.fir 295099:6]
  wire [9:0] _wrap_value_T_7 = rxBaudCount + 10'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 295101:6]
  wire  rxBaudWrap = txfifo_io_enq_ready & wrap_wrap_3; // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295098:4 Counter.scala 118:24 chipyard.TestHarness.RocketConfig.fir 295106:6 chipyard.TestHarness.RocketConfig.fir 295097:4]
  wire  _T_14 = rxState == 2'h2; // @[UARTAdapter.scala 83:49 chipyard.TestHarness.RocketConfig.fir 295108:4]
  wire  _T_15 = _T_14 & txfifo_io_enq_ready; // @[UARTAdapter.scala 83:61 chipyard.TestHarness.RocketConfig.fir 295109:4]
  wire  _T_16 = _T_15 & rxBaudWrap; // @[UARTAdapter.scala 83:84 chipyard.TestHarness.RocketConfig.fir 295110:4]
  reg [2:0] rxDataIdx; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295111:4]
  wire  wrap_wrap_4 = rxDataIdx == 3'h7; // @[Counter.scala 72:24 chipyard.TestHarness.RocketConfig.fir 295115:6]
  wire [2:0] _wrap_value_T_9 = rxDataIdx + 3'h1; // @[Counter.scala 76:24 chipyard.TestHarness.RocketConfig.fir 295117:6]
  wire  rxDataWrap = _T_16 & wrap_wrap_4; // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295114:4 Counter.scala 118:24 chipyard.TestHarness.RocketConfig.fir 295119:6 chipyard.TestHarness.RocketConfig.fir 295113:4]
  wire  _T_17 = 2'h0 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.RocketConfig.fir 295122:4]
  wire  _T_18 = rxBaudWrap & rxfifo_io_deq_valid; // @[UARTAdapter.scala 89:24 chipyard.TestHarness.RocketConfig.fir 295125:6]
  wire  _T_19 = 2'h1 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.RocketConfig.fir 295131:6]
  wire  _T_20 = 2'h2 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.RocketConfig.fir 295139:8]
  wire [7:0] _io_uart_rxd_T = rxfifo_io_deq_bits >> rxDataIdx; // @[UARTAdapter.scala 100:42 chipyard.TestHarness.RocketConfig.fir 295141:10]
  wire  _T_21 = rxDataWrap & rxBaudWrap; // @[UARTAdapter.scala 101:23 chipyard.TestHarness.RocketConfig.fir 295144:10]
  wire [1:0] _GEN_28 = _T_21 ? 2'h0 : rxState; // @[UARTAdapter.scala 101:38 chipyard.TestHarness.RocketConfig.fir 295145:10 UARTAdapter.scala 102:17 chipyard.TestHarness.RocketConfig.fir 295146:12 UARTAdapter.scala 79:24 chipyard.TestHarness.RocketConfig.fir 295094:4]
  wire  _GEN_29 = _T_20 ? _io_uart_rxd_T[0] : 1'h1; // @[Conditional.scala 39:67 chipyard.TestHarness.RocketConfig.fir 295140:8 UARTAdapter.scala 100:19 chipyard.TestHarness.RocketConfig.fir 295143:10 UARTAdapter.scala 85:15 chipyard.TestHarness.RocketConfig.fir 295121:4]
  wire  _GEN_31 = _T_19 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67 chipyard.TestHarness.RocketConfig.fir 295132:6 UARTAdapter.scala 94:19 chipyard.TestHarness.RocketConfig.fir 295133:8]
  wire  _rxfifo_io_deq_ready_T_1 = _T_14 & rxDataWrap; // @[UARTAdapter.scala 106:48 chipyard.TestHarness.RocketConfig.fir 295150:4]
  wire  _rxfifo_io_deq_ready_T_2 = _rxfifo_io_deq_ready_T_1 & rxBaudWrap; // @[UARTAdapter.scala 106:62 chipyard.TestHarness.RocketConfig.fir 295151:4]
  Queue_44_inTestHarness txfifo ( // @[UARTAdapter.scala 32:22 chipyard.TestHarness.RocketConfig.fir 295002:4]
    .clock(txfifo_clock),
    .reset(txfifo_reset),
    .io_enq_ready(txfifo_io_enq_ready),
    .io_enq_valid(txfifo_io_enq_valid),
    .io_enq_bits(txfifo_io_enq_bits),
    .io_deq_ready(txfifo_io_deq_ready),
    .io_deq_valid(txfifo_io_deq_valid),
    .io_deq_bits(txfifo_io_deq_bits)
  );
  Queue_44_inTestHarness rxfifo ( // @[UARTAdapter.scala 33:22 chipyard.TestHarness.RocketConfig.fir 295005:4]
    .clock(rxfifo_clock),
    .reset(rxfifo_reset),
    .io_enq_ready(rxfifo_io_enq_ready),
    .io_enq_valid(rxfifo_io_enq_valid),
    .io_enq_bits(rxfifo_io_enq_bits),
    .io_deq_ready(rxfifo_io_deq_ready),
    .io_deq_valid(rxfifo_io_deq_valid),
    .io_deq_bits(rxfifo_io_deq_bits)
  );
  SimUART #(.UARTNO(0)) sim ( // @[UARTAdapter.scala 108:19 chipyard.TestHarness.RocketConfig.fir 295154:4]
    .clock(sim_clock),
    .reset(sim_reset),
    .serial_in_ready(sim_serial_in_ready),
    .serial_in_valid(sim_serial_in_valid),
    .serial_in_bits(sim_serial_in_bits),
    .serial_out_ready(sim_serial_out_ready),
    .serial_out_valid(sim_serial_out_valid),
    .serial_out_bits(sim_serial_out_bits)
  );
  assign io_uart_rxd = _T_17 | _GEN_31; // @[Conditional.scala 40:58 chipyard.TestHarness.RocketConfig.fir 295123:4 UARTAdapter.scala 88:19 chipyard.TestHarness.RocketConfig.fir 295124:6]
  assign txfifo_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 295003:4]
  assign txfifo_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 295004:4]
  assign txfifo_io_enq_valid = _T_1 & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295015:4 Counter.scala 118:24 chipyard.TestHarness.RocketConfig.fir 295020:6 chipyard.TestHarness.RocketConfig.fir 295014:4]
  assign txfifo_io_enq_bits = txData; // @[UARTAdapter.scala 75:23 chipyard.TestHarness.RocketConfig.fir 295092:4]
  assign txfifo_io_deq_ready = sim_serial_out_ready; // @[UARTAdapter.scala 115:23 chipyard.TestHarness.RocketConfig.fir 295163:4]
  assign rxfifo_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 295006:4]
  assign rxfifo_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 295007:4]
  assign rxfifo_io_enq_valid = sim_serial_in_valid; // @[UARTAdapter.scala 118:23 chipyard.TestHarness.RocketConfig.fir 295165:4]
  assign rxfifo_io_enq_bits = sim_serial_in_bits; // @[UARTAdapter.scala 117:22 chipyard.TestHarness.RocketConfig.fir 295164:4]
  assign rxfifo_io_deq_ready = _rxfifo_io_deq_ready_T_2 & txfifo_io_enq_ready; // @[UARTAdapter.scala 106:76 chipyard.TestHarness.RocketConfig.fir 295152:4]
  assign sim_clock = clock; // @[UARTAdapter.scala 110:16 chipyard.TestHarness.RocketConfig.fir 295158:4]
  assign sim_reset = reset; // @[UARTAdapter.scala 111:25 chipyard.TestHarness.RocketConfig.fir 295159:4]
  assign sim_serial_in_ready = rxfifo_io_enq_ready; // @[UARTAdapter.scala 119:26 chipyard.TestHarness.RocketConfig.fir 295166:4]
  assign sim_serial_out_valid = txfifo_io_deq_valid; // @[UARTAdapter.scala 114:27 chipyard.TestHarness.RocketConfig.fir 295162:4]
  assign sim_serial_out_bits = txfifo_io_deq_bits; // @[UARTAdapter.scala 113:26 chipyard.TestHarness.RocketConfig.fir 295161:4]
  always @(posedge clock) begin
    if (reset) begin // @[UARTAdapter.scala 38:24 chipyard.TestHarness.RocketConfig.fir 295008:4]
      txState <= 2'h0; // @[UARTAdapter.scala 38:24 chipyard.TestHarness.RocketConfig.fir 295008:4]
    end else if (_T_8) begin // @[Conditional.scala 40:58 chipyard.TestHarness.RocketConfig.fir 295052:4]
      if (txSlackWrap) begin // @[UARTAdapter.scala 48:25 chipyard.TestHarness.RocketConfig.fir 295053:6]
        txState <= 2'h1; // @[UARTAdapter.scala 50:17 chipyard.TestHarness.RocketConfig.fir 295055:8]
      end
    end else if (_T_9) begin // @[Conditional.scala 39:67 chipyard.TestHarness.RocketConfig.fir 295060:6]
      if (txBaudWrap) begin // @[UARTAdapter.scala 54:24 chipyard.TestHarness.RocketConfig.fir 295061:8]
        txState <= 2'h2; // @[UARTAdapter.scala 55:17 chipyard.TestHarness.RocketConfig.fir 295062:10]
      end
    end else if (_T_10) begin // @[Conditional.scala 39:67 chipyard.TestHarness.RocketConfig.fir 295067:8]
      txState <= _GEN_12;
    end else begin
      txState <= _GEN_14;
    end
    if (_T_8) begin // @[Conditional.scala 40:58 chipyard.TestHarness.RocketConfig.fir 295052:4]
      if (txSlackWrap) begin // @[UARTAdapter.scala 48:25 chipyard.TestHarness.RocketConfig.fir 295053:6]
        txData <= 8'h0; // @[UARTAdapter.scala 49:17 chipyard.TestHarness.RocketConfig.fir 295054:8]
      end
    end else if (!(_T_9)) begin // @[Conditional.scala 39:67 chipyard.TestHarness.RocketConfig.fir 295060:6]
      if (_T_10) begin // @[Conditional.scala 39:67 chipyard.TestHarness.RocketConfig.fir 295067:8]
        if (txfifo_io_enq_ready) begin // @[UARTAdapter.scala 59:34 chipyard.TestHarness.RocketConfig.fir 295068:10]
          txData <= _txData_T_1; // @[UARTAdapter.scala 60:16 chipyard.TestHarness.RocketConfig.fir 295071:12]
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295012:4]
      txDataIdx <= 3'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295012:4]
    end else if (_T_1) begin // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295015:4]
      txDataIdx <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 295019:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295024:4]
      txBaudCount <= 10'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295024:4]
    end else if (_T_3) begin // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295027:4]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20 chipyard.TestHarness.RocketConfig.fir 295032:6]
        txBaudCount <= 10'h0; // @[Counter.scala 86:28 chipyard.TestHarness.RocketConfig.fir 295033:8]
      end else begin
        txBaudCount <= _wrap_value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 295031:6]
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295041:4]
      txSlackCount <= 2'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295041:4]
    end else if (_T_7) begin // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295044:4]
      txSlackCount <= _wrap_value_T_5; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 295048:6]
    end
    if (reset) begin // @[UARTAdapter.scala 79:24 chipyard.TestHarness.RocketConfig.fir 295094:4]
      rxState <= 2'h0; // @[UARTAdapter.scala 79:24 chipyard.TestHarness.RocketConfig.fir 295094:4]
    end else if (_T_17) begin // @[Conditional.scala 40:58 chipyard.TestHarness.RocketConfig.fir 295123:4]
      if (_T_18) begin // @[UARTAdapter.scala 89:48 chipyard.TestHarness.RocketConfig.fir 295126:6]
        rxState <= 2'h1; // @[UARTAdapter.scala 90:17 chipyard.TestHarness.RocketConfig.fir 295127:8]
      end
    end else if (_T_19) begin // @[Conditional.scala 39:67 chipyard.TestHarness.RocketConfig.fir 295132:6]
      if (rxBaudWrap) begin // @[UARTAdapter.scala 95:24 chipyard.TestHarness.RocketConfig.fir 295134:8]
        rxState <= 2'h2; // @[UARTAdapter.scala 96:17 chipyard.TestHarness.RocketConfig.fir 295135:10]
      end
    end else if (_T_20) begin // @[Conditional.scala 39:67 chipyard.TestHarness.RocketConfig.fir 295140:8]
      rxState <= _GEN_28;
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295095:4]
      rxBaudCount <= 10'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295095:4]
    end else if (txfifo_io_enq_ready) begin // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295098:4]
      if (wrap_wrap_3) begin // @[Counter.scala 86:20 chipyard.TestHarness.RocketConfig.fir 295103:6]
        rxBaudCount <= 10'h0; // @[Counter.scala 86:28 chipyard.TestHarness.RocketConfig.fir 295104:8]
      end else begin
        rxBaudCount <= _wrap_value_T_7; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 295102:6]
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295111:4]
      rxDataIdx <= 3'h0; // @[Counter.scala 60:40 chipyard.TestHarness.RocketConfig.fir 295111:4]
    end else if (_T_16) begin // @[Counter.scala 118:17 chipyard.TestHarness.RocketConfig.fir 295114:4]
      rxDataIdx <= _wrap_value_T_9; // @[Counter.scala 76:15 chipyard.TestHarness.RocketConfig.fir 295118:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  txState = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  txData = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  txDataIdx = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  txBaudCount = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  txSlackCount = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  rxState = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  rxBaudCount = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  rxDataIdx = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TestHarness( // @[chipyard.TestHarness.RocketConfig.fir 295168:2]
  input   clock, // @[chipyard.TestHarness.RocketConfig.fir 295169:4]
  input   reset, // @[chipyard.TestHarness.RocketConfig.fir 295170:4]
  output  io_success // @[chipyard.TestHarness.RocketConfig.fir 295171:4]
);
  wire  chiptop_jtag_TCK; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_jtag_TMS; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_jtag_TDI; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_jtag_TDO_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_jtag_TDO_driven; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_serial_tl_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_serial_tl_bits_in_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_serial_tl_bits_in_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [3:0] chiptop_serial_tl_bits_in_bits; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_serial_tl_bits_out_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_serial_tl_bits_out_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [3:0] chiptop_serial_tl_bits_out_bits; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_reset; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_aw_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_aw_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [3:0] chiptop_axi4_mem_0_bits_aw_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [31:0] chiptop_axi4_mem_0_bits_aw_bits_addr; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [7:0] chiptop_axi4_mem_0_bits_aw_bits_len; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [2:0] chiptop_axi4_mem_0_bits_aw_bits_size; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [1:0] chiptop_axi4_mem_0_bits_aw_bits_burst; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_aw_bits_lock; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [3:0] chiptop_axi4_mem_0_bits_aw_bits_cache; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [2:0] chiptop_axi4_mem_0_bits_aw_bits_prot; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [3:0] chiptop_axi4_mem_0_bits_aw_bits_qos; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_w_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_w_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [63:0] chiptop_axi4_mem_0_bits_w_bits_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [7:0] chiptop_axi4_mem_0_bits_w_bits_strb; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_w_bits_last; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_b_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_b_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [3:0] chiptop_axi4_mem_0_bits_b_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [1:0] chiptop_axi4_mem_0_bits_b_bits_resp; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_ar_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_ar_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [3:0] chiptop_axi4_mem_0_bits_ar_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [31:0] chiptop_axi4_mem_0_bits_ar_bits_addr; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [7:0] chiptop_axi4_mem_0_bits_ar_bits_len; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [2:0] chiptop_axi4_mem_0_bits_ar_bits_size; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [1:0] chiptop_axi4_mem_0_bits_ar_bits_burst; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_ar_bits_lock; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [3:0] chiptop_axi4_mem_0_bits_ar_bits_cache; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [2:0] chiptop_axi4_mem_0_bits_ar_bits_prot; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [3:0] chiptop_axi4_mem_0_bits_ar_bits_qos; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_r_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_r_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [3:0] chiptop_axi4_mem_0_bits_r_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [63:0] chiptop_axi4_mem_0_bits_r_bits_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire [1:0] chiptop_axi4_mem_0_bits_r_bits_resp; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_axi4_mem_0_bits_r_bits_last; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_uart_0_txd; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_uart_0_rxd; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_reset_wire_reset; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  chiptop_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
  wire  SimJTAG_clock; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire  SimJTAG_reset; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire  SimJTAG_jtag_TRSTn; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire  SimJTAG_jtag_TCK; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire  SimJTAG_jtag_TMS; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire  SimJTAG_jtag_TDI; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire  SimJTAG_jtag_TDO_data; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire  SimJTAG_jtag_TDO_driven; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire  SimJTAG_enable; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire  SimJTAG_init_done; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire [31:0] SimJTAG_exit; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 295202:4]
  wire  ram_clock; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire  ram_reset; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire  ram_io_ser_in_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire  ram_io_ser_in_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire [3:0] ram_io_ser_in_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire  ram_io_ser_out_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire  ram_io_ser_out_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire [3:0] ram_io_ser_out_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire  ram_io_tsi_ser_in_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire  ram_io_tsi_ser_in_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire [31:0] ram_io_tsi_ser_in_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire  ram_io_tsi_ser_out_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire  ram_io_tsi_ser_out_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire [31:0] ram_io_tsi_ser_out_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
  wire  success_sim_clock; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.RocketConfig.fir 295232:4]
  wire  success_sim_reset; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.RocketConfig.fir 295232:4]
  wire  success_sim_serial_in_ready; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.RocketConfig.fir 295232:4]
  wire  success_sim_serial_in_valid; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.RocketConfig.fir 295232:4]
  wire [31:0] success_sim_serial_in_bits; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.RocketConfig.fir 295232:4]
  wire  success_sim_serial_out_ready; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.RocketConfig.fir 295232:4]
  wire  success_sim_serial_out_valid; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.RocketConfig.fir 295232:4]
  wire [31:0] success_sim_serial_out_bits; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.RocketConfig.fir 295232:4]
  wire  success_sim_exit; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.RocketConfig.fir 295232:4]
  wire  simdram_clock; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_reset; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_aw_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_aw_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [3:0] simdram_axi_aw_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [31:0] simdram_axi_aw_bits_addr; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [7:0] simdram_axi_aw_bits_len; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [2:0] simdram_axi_aw_bits_size; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [1:0] simdram_axi_aw_bits_burst; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_aw_bits_lock; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [3:0] simdram_axi_aw_bits_cache; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [2:0] simdram_axi_aw_bits_prot; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [3:0] simdram_axi_aw_bits_qos; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_w_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_w_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [63:0] simdram_axi_w_bits_data; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [7:0] simdram_axi_w_bits_strb; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_w_bits_last; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_b_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_b_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [3:0] simdram_axi_b_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [1:0] simdram_axi_b_bits_resp; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_ar_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_ar_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [3:0] simdram_axi_ar_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [31:0] simdram_axi_ar_bits_addr; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [7:0] simdram_axi_ar_bits_len; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [2:0] simdram_axi_ar_bits_size; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [1:0] simdram_axi_ar_bits_burst; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_ar_bits_lock; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [3:0] simdram_axi_ar_bits_cache; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [2:0] simdram_axi_ar_bits_prot; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [3:0] simdram_axi_ar_bits_qos; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_r_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_r_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [3:0] simdram_axi_r_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [63:0] simdram_axi_r_bits_data; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire [1:0] simdram_axi_r_bits_resp; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  simdram_axi_r_bits_last; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
  wire  uart_sim_0_clock; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.RocketConfig.fir 295255:4]
  wire  uart_sim_0_reset; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.RocketConfig.fir 295255:4]
  wire  uart_sim_0_io_uart_txd; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.RocketConfig.fir 295255:4]
  wire  uart_sim_0_io_uart_rxd; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.RocketConfig.fir 295255:4]
  wire  dtm_success = SimJTAG_exit == 32'h1; // @[Periphery.scala 233:26 chipyard.TestHarness.RocketConfig.fir 295206:4]
  wire  _T_2 = ~reset; // @[HarnessBinders.scala 190:105 chipyard.TestHarness.RocketConfig.fir 295194:4]
  wire  _T_3 = SimJTAG_exit >= 32'h2; // @[Periphery.scala 234:19 chipyard.TestHarness.RocketConfig.fir 295208:4]
  wire [31:0] _T_4 = {{1'd0}, SimJTAG_exit[31:1]}; // @[Periphery.scala 235:59 chipyard.TestHarness.RocketConfig.fir 295210:6]
  ChipTop chiptop ( // @[TestHarness.scala 34:19 chipyard.TestHarness.RocketConfig.fir 295173:4]
    .jtag_TCK(chiptop_jtag_TCK),
    .jtag_TMS(chiptop_jtag_TMS),
    .jtag_TDI(chiptop_jtag_TDI),
    .jtag_TDO_data(chiptop_jtag_TDO_data),
    .jtag_TDO_driven(chiptop_jtag_TDO_driven),
    .serial_tl_clock(chiptop_serial_tl_clock),
    .serial_tl_bits_in_ready(chiptop_serial_tl_bits_in_ready),
    .serial_tl_bits_in_valid(chiptop_serial_tl_bits_in_valid),
    .serial_tl_bits_in_bits(chiptop_serial_tl_bits_in_bits),
    .serial_tl_bits_out_ready(chiptop_serial_tl_bits_out_ready),
    .serial_tl_bits_out_valid(chiptop_serial_tl_bits_out_valid),
    .serial_tl_bits_out_bits(chiptop_serial_tl_bits_out_bits),
    .axi4_mem_0_clock(chiptop_axi4_mem_0_clock),
    .axi4_mem_0_reset(chiptop_axi4_mem_0_reset),
    .axi4_mem_0_bits_aw_ready(chiptop_axi4_mem_0_bits_aw_ready),
    .axi4_mem_0_bits_aw_valid(chiptop_axi4_mem_0_bits_aw_valid),
    .axi4_mem_0_bits_aw_bits_id(chiptop_axi4_mem_0_bits_aw_bits_id),
    .axi4_mem_0_bits_aw_bits_addr(chiptop_axi4_mem_0_bits_aw_bits_addr),
    .axi4_mem_0_bits_aw_bits_len(chiptop_axi4_mem_0_bits_aw_bits_len),
    .axi4_mem_0_bits_aw_bits_size(chiptop_axi4_mem_0_bits_aw_bits_size),
    .axi4_mem_0_bits_aw_bits_burst(chiptop_axi4_mem_0_bits_aw_bits_burst),
    .axi4_mem_0_bits_aw_bits_lock(chiptop_axi4_mem_0_bits_aw_bits_lock),
    .axi4_mem_0_bits_aw_bits_cache(chiptop_axi4_mem_0_bits_aw_bits_cache),
    .axi4_mem_0_bits_aw_bits_prot(chiptop_axi4_mem_0_bits_aw_bits_prot),
    .axi4_mem_0_bits_aw_bits_qos(chiptop_axi4_mem_0_bits_aw_bits_qos),
    .axi4_mem_0_bits_w_ready(chiptop_axi4_mem_0_bits_w_ready),
    .axi4_mem_0_bits_w_valid(chiptop_axi4_mem_0_bits_w_valid),
    .axi4_mem_0_bits_w_bits_data(chiptop_axi4_mem_0_bits_w_bits_data),
    .axi4_mem_0_bits_w_bits_strb(chiptop_axi4_mem_0_bits_w_bits_strb),
    .axi4_mem_0_bits_w_bits_last(chiptop_axi4_mem_0_bits_w_bits_last),
    .axi4_mem_0_bits_b_ready(chiptop_axi4_mem_0_bits_b_ready),
    .axi4_mem_0_bits_b_valid(chiptop_axi4_mem_0_bits_b_valid),
    .axi4_mem_0_bits_b_bits_id(chiptop_axi4_mem_0_bits_b_bits_id),
    .axi4_mem_0_bits_b_bits_resp(chiptop_axi4_mem_0_bits_b_bits_resp),
    .axi4_mem_0_bits_ar_ready(chiptop_axi4_mem_0_bits_ar_ready),
    .axi4_mem_0_bits_ar_valid(chiptop_axi4_mem_0_bits_ar_valid),
    .axi4_mem_0_bits_ar_bits_id(chiptop_axi4_mem_0_bits_ar_bits_id),
    .axi4_mem_0_bits_ar_bits_addr(chiptop_axi4_mem_0_bits_ar_bits_addr),
    .axi4_mem_0_bits_ar_bits_len(chiptop_axi4_mem_0_bits_ar_bits_len),
    .axi4_mem_0_bits_ar_bits_size(chiptop_axi4_mem_0_bits_ar_bits_size),
    .axi4_mem_0_bits_ar_bits_burst(chiptop_axi4_mem_0_bits_ar_bits_burst),
    .axi4_mem_0_bits_ar_bits_lock(chiptop_axi4_mem_0_bits_ar_bits_lock),
    .axi4_mem_0_bits_ar_bits_cache(chiptop_axi4_mem_0_bits_ar_bits_cache),
    .axi4_mem_0_bits_ar_bits_prot(chiptop_axi4_mem_0_bits_ar_bits_prot),
    .axi4_mem_0_bits_ar_bits_qos(chiptop_axi4_mem_0_bits_ar_bits_qos),
    .axi4_mem_0_bits_r_ready(chiptop_axi4_mem_0_bits_r_ready),
    .axi4_mem_0_bits_r_valid(chiptop_axi4_mem_0_bits_r_valid),
    .axi4_mem_0_bits_r_bits_id(chiptop_axi4_mem_0_bits_r_bits_id),
    .axi4_mem_0_bits_r_bits_data(chiptop_axi4_mem_0_bits_r_bits_data),
    .axi4_mem_0_bits_r_bits_resp(chiptop_axi4_mem_0_bits_r_bits_resp),
    .axi4_mem_0_bits_r_bits_last(chiptop_axi4_mem_0_bits_r_bits_last),
    .uart_0_txd(chiptop_uart_0_txd),
    .uart_0_rxd(chiptop_uart_0_rxd),
    .reset_wire_reset(chiptop_reset_wire_reset),
    .clock(chiptop_clock)
  );
  SimJTAG #(.TICK_DELAY(3)) SimJTAG ( // @[HarnessBinders.scala 190:26 chipyard.TestHarness.RocketConfig.fir 295185:4]
    .clock(SimJTAG_clock),
    .reset(SimJTAG_reset),
    .jtag_TRSTn(SimJTAG_jtag_TRSTn),
    .jtag_TCK(SimJTAG_jtag_TCK),
    .jtag_TMS(SimJTAG_jtag_TMS),
    .jtag_TDI(SimJTAG_jtag_TDI),
    .jtag_TDO_data(SimJTAG_jtag_TDO_data),
    .jtag_TDO_driven(SimJTAG_jtag_TDO_driven),
    .enable(SimJTAG_enable),
    .init_done(SimJTAG_init_done),
    .exit(SimJTAG_exit)
  );
  plusarg_reader #(.FORMAT("jtag_rbb_enable=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.RocketConfig.fir 295202:4]
    .out(plusarg_reader_out)
  );
  SerialRAM_inTestHarness ram ( // @[SerialAdapter.scala 27:26 chipyard.TestHarness.RocketConfig.fir 295222:4]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_ser_in_ready(ram_io_ser_in_ready),
    .io_ser_in_valid(ram_io_ser_in_valid),
    .io_ser_in_bits(ram_io_ser_in_bits),
    .io_ser_out_ready(ram_io_ser_out_ready),
    .io_ser_out_valid(ram_io_ser_out_valid),
    .io_ser_out_bits(ram_io_ser_out_bits),
    .io_tsi_ser_in_ready(ram_io_tsi_ser_in_ready),
    .io_tsi_ser_in_valid(ram_io_tsi_ser_in_valid),
    .io_tsi_ser_in_bits(ram_io_tsi_ser_in_bits),
    .io_tsi_ser_out_ready(ram_io_tsi_ser_out_ready),
    .io_tsi_ser_out_valid(ram_io_tsi_ser_out_valid),
    .io_tsi_ser_out_bits(ram_io_tsi_ser_out_bits)
  );
  SimSerial success_sim ( // @[SerialAdapter.scala 37:23 chipyard.TestHarness.RocketConfig.fir 295232:4]
    .clock(success_sim_clock),
    .reset(success_sim_reset),
    .serial_in_ready(success_sim_serial_in_ready),
    .serial_in_valid(success_sim_serial_in_valid),
    .serial_in_bits(success_sim_serial_in_bits),
    .serial_out_ready(success_sim_serial_out_ready),
    .serial_out_valid(success_sim_serial_out_valid),
    .serial_out_bits(success_sim_serial_out_bits),
    .exit(success_sim_exit)
  );
  SimDRAM #(.LINE_SIZE(64), .ID_BITS(4), .ADDR_BITS(32), .MEM_SIZE(268435456), .DATA_BITS(64)) simdram ( // @[HarnessBinders.scala 146:23 chipyard.TestHarness.RocketConfig.fir 295248:4]
    .clock(simdram_clock),
    .reset(simdram_reset),
    .axi_aw_ready(simdram_axi_aw_ready),
    .axi_aw_valid(simdram_axi_aw_valid),
    .axi_aw_bits_id(simdram_axi_aw_bits_id),
    .axi_aw_bits_addr(simdram_axi_aw_bits_addr),
    .axi_aw_bits_len(simdram_axi_aw_bits_len),
    .axi_aw_bits_size(simdram_axi_aw_bits_size),
    .axi_aw_bits_burst(simdram_axi_aw_bits_burst),
    .axi_aw_bits_lock(simdram_axi_aw_bits_lock),
    .axi_aw_bits_cache(simdram_axi_aw_bits_cache),
    .axi_aw_bits_prot(simdram_axi_aw_bits_prot),
    .axi_aw_bits_qos(simdram_axi_aw_bits_qos),
    .axi_w_ready(simdram_axi_w_ready),
    .axi_w_valid(simdram_axi_w_valid),
    .axi_w_bits_data(simdram_axi_w_bits_data),
    .axi_w_bits_strb(simdram_axi_w_bits_strb),
    .axi_w_bits_last(simdram_axi_w_bits_last),
    .axi_b_ready(simdram_axi_b_ready),
    .axi_b_valid(simdram_axi_b_valid),
    .axi_b_bits_id(simdram_axi_b_bits_id),
    .axi_b_bits_resp(simdram_axi_b_bits_resp),
    .axi_ar_ready(simdram_axi_ar_ready),
    .axi_ar_valid(simdram_axi_ar_valid),
    .axi_ar_bits_id(simdram_axi_ar_bits_id),
    .axi_ar_bits_addr(simdram_axi_ar_bits_addr),
    .axi_ar_bits_len(simdram_axi_ar_bits_len),
    .axi_ar_bits_size(simdram_axi_ar_bits_size),
    .axi_ar_bits_burst(simdram_axi_ar_bits_burst),
    .axi_ar_bits_lock(simdram_axi_ar_bits_lock),
    .axi_ar_bits_cache(simdram_axi_ar_bits_cache),
    .axi_ar_bits_prot(simdram_axi_ar_bits_prot),
    .axi_ar_bits_qos(simdram_axi_ar_bits_qos),
    .axi_r_ready(simdram_axi_r_ready),
    .axi_r_valid(simdram_axi_r_valid),
    .axi_r_bits_id(simdram_axi_r_bits_id),
    .axi_r_bits_data(simdram_axi_r_bits_data),
    .axi_r_bits_resp(simdram_axi_r_bits_resp),
    .axi_r_bits_last(simdram_axi_r_bits_last)
  );
  UARTAdapter_inTestHarness uart_sim_0 ( // @[UARTAdapter.scala 132:28 chipyard.TestHarness.RocketConfig.fir 295255:4]
    .clock(uart_sim_0_clock),
    .reset(uart_sim_0_reset),
    .io_uart_txd(uart_sim_0_io_uart_txd),
    .io_uart_rxd(uart_sim_0_io_uart_rxd)
  );
  assign io_success = success_sim_exit | dtm_success; // @[HarnessBinders.scala 236:22 chipyard.TestHarness.RocketConfig.fir 295245:4 HarnessBinders.scala 236:35 chipyard.TestHarness.RocketConfig.fir 295246:6]
  assign chiptop_jtag_TCK = SimJTAG_jtag_TCK; // @[Periphery.scala 220:15 chipyard.TestHarness.RocketConfig.fir 295195:4]
  assign chiptop_jtag_TMS = SimJTAG_jtag_TMS; // @[Periphery.scala 221:15 chipyard.TestHarness.RocketConfig.fir 295196:4]
  assign chiptop_jtag_TDI = SimJTAG_jtag_TDI; // @[Periphery.scala 222:15 chipyard.TestHarness.RocketConfig.fir 295197:4]
  assign chiptop_serial_tl_bits_in_valid = ram_io_ser_in_valid; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.RocketConfig.fir 295229:4]
  assign chiptop_serial_tl_bits_in_bits = ram_io_ser_in_bits; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.RocketConfig.fir 295228:4]
  assign chiptop_serial_tl_bits_out_ready = ram_io_ser_out_ready; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.RocketConfig.fir 295227:4]
  assign chiptop_axi4_mem_0_bits_aw_ready = simdram_axi_aw_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_axi4_mem_0_bits_w_ready = simdram_axi_w_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_axi4_mem_0_bits_b_valid = simdram_axi_b_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_axi4_mem_0_bits_b_bits_id = simdram_axi_b_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_axi4_mem_0_bits_b_bits_resp = simdram_axi_b_bits_resp; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_axi4_mem_0_bits_ar_ready = simdram_axi_ar_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_axi4_mem_0_bits_r_valid = simdram_axi_r_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_axi4_mem_0_bits_r_bits_id = simdram_axi_r_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_axi4_mem_0_bits_r_bits_data = simdram_axi_r_bits_data; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_axi4_mem_0_bits_r_bits_resp = simdram_axi_r_bits_resp; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_axi4_mem_0_bits_r_bits_last = simdram_axi_r_bits_last; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign chiptop_uart_0_rxd = uart_sim_0_io_uart_rxd; // @[UARTAdapter.scala 135:18 chipyard.TestHarness.RocketConfig.fir 295259:4]
  assign chiptop_reset_wire_reset = reset; // @[TestHarness.scala 41:24 chipyard.TestHarness.RocketConfig.fir 295177:4]
  assign chiptop_clock = clock; // @[Clocks.scala 106:18 chipyard.TestHarness.RocketConfig.fir 295179:4]
  assign SimJTAG_clock = clock; // @[Periphery.scala 225:14 chipyard.TestHarness.RocketConfig.fir 295200:4]
  assign SimJTAG_reset = reset; // @[HarnessBinders.scala 190:97 chipyard.TestHarness.RocketConfig.fir 295192:4]
  assign SimJTAG_jtag_TDO_data = chiptop_jtag_TDO_data; // @[Periphery.scala 223:17 chipyard.TestHarness.RocketConfig.fir 295199:4]
  assign SimJTAG_jtag_TDO_driven = chiptop_jtag_TDO_driven; // @[Periphery.scala 223:17 chipyard.TestHarness.RocketConfig.fir 295198:4]
  assign SimJTAG_enable = plusarg_reader_out[0]; // @[Periphery.scala 228:18 chipyard.TestHarness.RocketConfig.fir 295204:4]
  assign SimJTAG_init_done = ~reset; // @[HarnessBinders.scala 190:105 chipyard.TestHarness.RocketConfig.fir 295194:4]
  assign ram_clock = chiptop_serial_tl_clock; // @[chipyard.TestHarness.RocketConfig.fir 295223:4]
  assign ram_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 295175:4 chipyard.TestHarness.RocketConfig.fir 295176:4]
  assign ram_io_ser_in_ready = chiptop_serial_tl_bits_in_ready; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.RocketConfig.fir 295230:4]
  assign ram_io_ser_out_valid = chiptop_serial_tl_bits_out_valid; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.RocketConfig.fir 295226:4]
  assign ram_io_ser_out_bits = chiptop_serial_tl_bits_out_bits; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.RocketConfig.fir 295225:4]
  assign ram_io_tsi_ser_in_valid = success_sim_serial_in_valid; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.RocketConfig.fir 295243:4]
  assign ram_io_tsi_ser_in_bits = success_sim_serial_in_bits; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.RocketConfig.fir 295242:4]
  assign ram_io_tsi_ser_out_ready = success_sim_serial_out_ready; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.RocketConfig.fir 295241:4]
  assign success_sim_clock = chiptop_serial_tl_clock; // @[SerialAdapter.scala 38:20 chipyard.TestHarness.RocketConfig.fir 295237:4]
  assign success_sim_reset = reset; // @[HarnessBinders.scala 235:103 chipyard.TestHarness.RocketConfig.fir 295231:4]
  assign success_sim_serial_in_ready = ram_io_tsi_ser_in_ready; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.RocketConfig.fir 295244:4]
  assign success_sim_serial_out_valid = ram_io_tsi_ser_out_valid; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.RocketConfig.fir 295240:4]
  assign success_sim_serial_out_bits = ram_io_tsi_ser_out_bits; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.RocketConfig.fir 295239:4]
  assign simdram_clock = chiptop_axi4_mem_0_clock; // @[HarnessBinders.scala 148:20 chipyard.TestHarness.RocketConfig.fir 295253:4]
  assign simdram_reset = chiptop_axi4_mem_0_reset; // @[HarnessBinders.scala 149:20 chipyard.TestHarness.RocketConfig.fir 295254:4]
  assign simdram_axi_aw_valid = chiptop_axi4_mem_0_bits_aw_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_aw_bits_id = chiptop_axi4_mem_0_bits_aw_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_aw_bits_addr = chiptop_axi4_mem_0_bits_aw_bits_addr; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_aw_bits_len = chiptop_axi4_mem_0_bits_aw_bits_len; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_aw_bits_size = chiptop_axi4_mem_0_bits_aw_bits_size; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_aw_bits_burst = chiptop_axi4_mem_0_bits_aw_bits_burst; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_aw_bits_lock = chiptop_axi4_mem_0_bits_aw_bits_lock; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_aw_bits_cache = chiptop_axi4_mem_0_bits_aw_bits_cache; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_aw_bits_prot = chiptop_axi4_mem_0_bits_aw_bits_prot; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_aw_bits_qos = chiptop_axi4_mem_0_bits_aw_bits_qos; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_w_valid = chiptop_axi4_mem_0_bits_w_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_w_bits_data = chiptop_axi4_mem_0_bits_w_bits_data; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_w_bits_strb = chiptop_axi4_mem_0_bits_w_bits_strb; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_w_bits_last = chiptop_axi4_mem_0_bits_w_bits_last; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_b_ready = chiptop_axi4_mem_0_bits_b_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_ar_valid = chiptop_axi4_mem_0_bits_ar_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_ar_bits_id = chiptop_axi4_mem_0_bits_ar_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_ar_bits_addr = chiptop_axi4_mem_0_bits_ar_bits_addr; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_ar_bits_len = chiptop_axi4_mem_0_bits_ar_bits_len; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_ar_bits_size = chiptop_axi4_mem_0_bits_ar_bits_size; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_ar_bits_burst = chiptop_axi4_mem_0_bits_ar_bits_burst; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_ar_bits_lock = chiptop_axi4_mem_0_bits_ar_bits_lock; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_ar_bits_cache = chiptop_axi4_mem_0_bits_ar_bits_cache; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_ar_bits_prot = chiptop_axi4_mem_0_bits_ar_bits_prot; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_ar_bits_qos = chiptop_axi4_mem_0_bits_ar_bits_qos; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign simdram_axi_r_ready = chiptop_axi4_mem_0_bits_r_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.RocketConfig.fir 295252:4]
  assign uart_sim_0_clock = clock; // @[chipyard.TestHarness.RocketConfig.fir 295256:4]
  assign uart_sim_0_reset = reset; // @[chipyard.TestHarness.RocketConfig.fir 295257:4]
  assign uart_sim_0_io_uart_txd = chiptop_uart_0_txd; // @[UARTAdapter.scala 134:28 chipyard.TestHarness.RocketConfig.fir 295258:4]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & _T_2) begin
          $fwrite(32'h80000002,"*** FAILED *** (exit code = %d)\n",_T_4); // @[Periphery.scala 235:13 chipyard.TestHarness.RocketConfig.fir 295214:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3 & _T_2) begin
          $fatal; // @[Periphery.scala 236:11 chipyard.TestHarness.RocketConfig.fir 295219:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module mem_inTestHarness(
  input  [8:0] RW0_addr,
  input        RW0_en,
  input        RW0_clk,
  input        RW0_wmode,
  input  [7:0] RW0_wdata_0,
  input  [7:0] RW0_wdata_1,
  input  [7:0] RW0_wdata_2,
  input  [7:0] RW0_wdata_3,
  input  [7:0] RW0_wdata_4,
  input  [7:0] RW0_wdata_5,
  input  [7:0] RW0_wdata_6,
  input  [7:0] RW0_wdata_7,
  output [7:0] RW0_rdata_0,
  output [7:0] RW0_rdata_1,
  output [7:0] RW0_rdata_2,
  output [7:0] RW0_rdata_3,
  output [7:0] RW0_rdata_4,
  output [7:0] RW0_rdata_5,
  output [7:0] RW0_rdata_6,
  output [7:0] RW0_rdata_7,
  input        RW0_wmask_0,
  input        RW0_wmask_1,
  input        RW0_wmask_2,
  input        RW0_wmask_3,
  input        RW0_wmask_4,
  input        RW0_wmask_5,
  input        RW0_wmask_6,
  input        RW0_wmask_7
);
  wire [8:0] mem_ext_RW0_addr;
  wire  mem_ext_RW0_en;
  wire  mem_ext_RW0_clk;
  wire  mem_ext_RW0_wmode;
  wire [63:0] mem_ext_RW0_wdata;
  wire [63:0] mem_ext_RW0_rdata;
  wire [7:0] mem_ext_RW0_wmask;
  wire [31:0] _GEN_4 = {RW0_wdata_7,RW0_wdata_6,RW0_wdata_5,RW0_wdata_4};
  wire [31:0] _GEN_5 = {RW0_wdata_3,RW0_wdata_2,RW0_wdata_1,RW0_wdata_0};
  wire [3:0] _GEN_10 = {RW0_wmask_7,RW0_wmask_6,RW0_wmask_5,RW0_wmask_4};
  wire [3:0] _GEN_11 = {RW0_wmask_3,RW0_wmask_2,RW0_wmask_1,RW0_wmask_0};
  mem_ext mem_ext (
    .RW0_addr(mem_ext_RW0_addr),
    .RW0_en(mem_ext_RW0_en),
    .RW0_clk(mem_ext_RW0_clk),
    .RW0_wmode(mem_ext_RW0_wmode),
    .RW0_wdata(mem_ext_RW0_wdata),
    .RW0_rdata(mem_ext_RW0_rdata),
    .RW0_wmask(mem_ext_RW0_wmask)
  );
  assign mem_ext_RW0_clk = RW0_clk;
  assign mem_ext_RW0_en = RW0_en;
  assign mem_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = mem_ext_RW0_rdata[7:0];
  assign RW0_rdata_1 = mem_ext_RW0_rdata[15:8];
  assign RW0_rdata_2 = mem_ext_RW0_rdata[23:16];
  assign RW0_rdata_3 = mem_ext_RW0_rdata[31:24];
  assign RW0_rdata_4 = mem_ext_RW0_rdata[39:32];
  assign RW0_rdata_5 = mem_ext_RW0_rdata[47:40];
  assign RW0_rdata_6 = mem_ext_RW0_rdata[55:48];
  assign RW0_rdata_7 = mem_ext_RW0_rdata[63:56];
  assign mem_ext_RW0_wmode = RW0_wmode;
  assign mem_ext_RW0_wdata = {_GEN_4,_GEN_5};
  assign mem_ext_RW0_wmask = {_GEN_10,_GEN_11};
endmodule
