module Queue_5_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 27698:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 27699:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 27700:4]
  output        io_enq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  input         io_enq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  input  [1:0]  io_enq_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  input  [6:0]  io_enq_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  input  [31:0] io_enq_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  input         io_deq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  output        io_deq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  output [1:0]  io_deq_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  output [1:0]  io_deq_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  output [6:0]  io_deq_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  output        io_deq_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  output        io_deq_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  output [31:0] io_deq_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 27701:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  reg [1:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  reg [6:0] ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire [6:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire [6:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  reg  ram_sink [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  reg [31:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 27704:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 27705:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 27706:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.TinyRocketConfig.fir 27707:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.TinyRocketConfig.fir 27708:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.TinyRocketConfig.fir 27709:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.TinyRocketConfig.fir 27710:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 27711:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 27714:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 27729:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 27735:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.TinyRocketConfig.fir 27738:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  assign ram_param_MPORT_data = 2'h0;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_addr = value_1;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  assign ram_sink_MPORT_data = 1'h0;
  assign ram_sink_MPORT_addr = value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  assign ram_denied_MPORT_data = 1'h0;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.TinyRocketConfig.fir 27744:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.TinyRocketConfig.fir 27742:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 27754:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 27753:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 27752:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 27751:4]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 27750:4]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 27749:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 27748:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 27747:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 27703:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 27704:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 27704:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.TinyRocketConfig.fir 27717:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 27730:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 27705:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 27705:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.TinyRocketConfig.fir 27732:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 27736:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 27706:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 27706:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.TinyRocketConfig.fir 27739:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.TinyRocketConfig.fir 27740:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_6_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 32859:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 32860:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 32861:4]
  output        io_enq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  input         io_enq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  input  [3:0]  io_enq_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  input  [31:0] io_enq_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  input  [3:0]  io_enq_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  input  [31:0] io_enq_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  input         io_deq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  output        io_deq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  output [3:0]  io_deq_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  output        io_deq_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  output [31:0] io_deq_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  output [3:0]  io_deq_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  output [31:0] io_deq_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 32862:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  reg  ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  reg [31:0] ram_address [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [31:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  reg [3:0] ram_mask [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [3:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [3:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  reg [31:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32865:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32866:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 32867:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.TinyRocketConfig.fir 32868:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.TinyRocketConfig.fir 32869:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.TinyRocketConfig.fir 32870:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.TinyRocketConfig.fir 32871:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 32872:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 32875:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 32890:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 32896:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.TinyRocketConfig.fir 32899:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  assign ram_param_MPORT_data = 3'h0;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  assign ram_source_MPORT_data = 1'h0;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.TinyRocketConfig.fir 32905:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.TinyRocketConfig.fir 32903:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32915:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32914:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32913:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32912:4]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32911:4]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32910:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32909:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32908:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32864:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32865:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32865:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.TinyRocketConfig.fir 32878:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 32891:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32866:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32866:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.TinyRocketConfig.fir 32893:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 32897:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 32867:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 32867:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.TinyRocketConfig.fir 32900:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.TinyRocketConfig.fir 32901:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_7_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 32923:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 32924:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 32925:4]
  output        io_enq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  input         io_enq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  input  [1:0]  io_enq_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  input  [3:0]  io_enq_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  input         io_enq_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  input         io_enq_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  input         io_enq_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  input  [31:0] io_enq_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  input         io_deq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  output        io_deq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  output [1:0]  io_deq_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  output [3:0]  io_deq_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  output        io_deq_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  output        io_deq_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  output        io_deq_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  output [31:0] io_deq_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 32926:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  reg  ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  reg  ram_sink [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  reg [31:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32929:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32930:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 32931:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.TinyRocketConfig.fir 32932:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.TinyRocketConfig.fir 32933:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.TinyRocketConfig.fir 32934:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.TinyRocketConfig.fir 32935:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 32936:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 32939:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 32954:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 32960:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.TinyRocketConfig.fir 32963:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_addr = value_1;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  assign ram_sink_MPORT_data = io_enq_bits_sink;
  assign ram_sink_MPORT_addr = value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.TinyRocketConfig.fir 32969:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.TinyRocketConfig.fir 32967:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32979:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32978:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32977:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32976:4]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32975:4]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32974:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32973:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 32972:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 32928:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32929:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32929:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.TinyRocketConfig.fir 32942:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 32955:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32930:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 32930:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.TinyRocketConfig.fir 32957:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 32961:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 32931:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 32931:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.TinyRocketConfig.fir 32964:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.TinyRocketConfig.fir 32965:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HellaPeekingArbiter_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 185005:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 185006:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 185007:4]
  output        io_in_1_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input         io_in_1_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [2:0]  io_in_1_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [2:0]  io_in_1_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [3:0]  io_in_1_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [1:0]  io_in_1_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [31:0] io_in_1_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input         io_in_1_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [3:0]  io_in_1_bits_union, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input         io_in_1_bits_last, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output        io_in_4_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input         io_in_4_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [2:0]  io_in_4_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [2:0]  io_in_4_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [3:0]  io_in_4_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [1:0]  io_in_4_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [31:0] io_in_4_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [31:0] io_in_4_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input         io_in_4_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input  [3:0]  io_in_4_bits_union, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input         io_in_4_bits_last, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  input         io_out_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output        io_out_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output [2:0]  io_out_bits_chanId, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output [2:0]  io_out_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output [2:0]  io_out_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output [3:0]  io_out_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output [1:0]  io_out_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output [31:0] io_out_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output [31:0] io_out_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output        io_out_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output [3:0]  io_out_bits_union, // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
  output        io_out_bits_last // @[chipyard.TestHarness.TinyRocketConfig.fir 185008:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lockIdx; // @[Arbiters.scala 25:20 chipyard.TestHarness.TinyRocketConfig.fir 185013:4]
  reg  locked; // @[Arbiters.scala 26:19 chipyard.TestHarness.TinyRocketConfig.fir 185014:4]
  wire [2:0] choice = io_in_1_valid ? 3'h1 : 3'h4; // @[Mux.scala 47:69 chipyard.TestHarness.TinyRocketConfig.fir 185017:4]
  wire [2:0] chosen = locked ? lockIdx : choice; // @[Arbiters.scala 36:19 chipyard.TestHarness.TinyRocketConfig.fir 185019:4]
  wire  _io_in_1_ready_T = chosen == 3'h1; // @[Arbiters.scala 39:46 chipyard.TestHarness.TinyRocketConfig.fir 185023:4]
  wire  _io_in_4_ready_T = chosen == 3'h4; // @[Arbiters.scala 39:46 chipyard.TestHarness.TinyRocketConfig.fir 185032:4]
  wire [2:0] _GEN_14 = 3'h1 == chosen ? 3'h3 : 3'h4; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [2:0] _GEN_15 = 3'h1 == chosen ? io_in_1_bits_opcode : 3'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [2:0] _GEN_16 = 3'h1 == chosen ? io_in_1_bits_param : 3'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [3:0] _GEN_17 = 3'h1 == chosen ? io_in_1_bits_size : 4'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [1:0] _GEN_18 = 3'h1 == chosen ? io_in_1_bits_source : 2'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [31:0] _GEN_20 = 3'h1 == chosen ? io_in_1_bits_data : 32'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [3:0] _GEN_22 = 3'h1 == chosen ? io_in_1_bits_union : 4'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire  _GEN_23 = 3'h1 == chosen ? io_in_1_bits_last : 1'h1; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire  _GEN_25 = 3'h2 == chosen ? 1'h0 : 3'h1 == chosen & io_in_1_valid; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [2:0] _GEN_26 = 3'h2 == chosen ? 3'h2 : _GEN_14; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [2:0] _GEN_27 = 3'h2 == chosen ? 3'h0 : _GEN_15; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [2:0] _GEN_28 = 3'h2 == chosen ? 3'h0 : _GEN_16; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [3:0] _GEN_29 = 3'h2 == chosen ? 4'h0 : _GEN_17; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [1:0] _GEN_30 = 3'h2 == chosen ? 2'h0 : _GEN_18; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [31:0] _GEN_32 = 3'h2 == chosen ? 32'h0 : _GEN_20; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire  _GEN_33 = 3'h2 == chosen ? 1'h0 : 3'h1 == chosen & io_in_1_bits_corrupt; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [3:0] _GEN_34 = 3'h2 == chosen ? 4'h0 : _GEN_22; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire  _GEN_37 = 3'h3 == chosen ? 1'h0 : _GEN_25; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [2:0] _GEN_38 = 3'h3 == chosen ? 3'h1 : _GEN_26; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [2:0] _GEN_39 = 3'h3 == chosen ? 3'h0 : _GEN_27; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [2:0] _GEN_40 = 3'h3 == chosen ? 3'h0 : _GEN_28; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [3:0] _GEN_41 = 3'h3 == chosen ? 4'h0 : _GEN_29; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [1:0] _GEN_42 = 3'h3 == chosen ? 2'h0 : _GEN_30; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [31:0] _GEN_44 = 3'h3 == chosen ? 32'h0 : _GEN_32; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire  _GEN_45 = 3'h3 == chosen ? 1'h0 : _GEN_33; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire [3:0] _GEN_46 = 3'h3 == chosen ? 4'h0 : _GEN_34; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 185037:4]
  wire  _T_1 = ~locked; // @[Arbiters.scala 59:11 chipyard.TestHarness.TinyRocketConfig.fir 185039:6]
  wire  _GEN_61 = _T_1 | locked; // @[Arbiters.scala 59:50 chipyard.TestHarness.TinyRocketConfig.fir 185041:6 Arbiters.scala 61:14 chipyard.TestHarness.TinyRocketConfig.fir 185043:8 Arbiters.scala 26:19 chipyard.TestHarness.TinyRocketConfig.fir 185014:4]
  assign io_in_1_ready = io_out_ready & _io_in_1_ready_T; // @[Arbiters.scala 39:36 chipyard.TestHarness.TinyRocketConfig.fir 185024:4]
  assign io_in_4_ready = io_out_ready & _io_in_4_ready_T; // @[Arbiters.scala 39:36 chipyard.TestHarness.TinyRocketConfig.fir 185033:4]
  assign io_out_valid = 3'h4 == chosen ? io_in_4_valid : _GEN_37; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  assign io_out_bits_chanId = 3'h4 == chosen ? 3'h0 : _GEN_38; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  assign io_out_bits_opcode = 3'h4 == chosen ? io_in_4_bits_opcode : _GEN_39; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  assign io_out_bits_param = 3'h4 == chosen ? io_in_4_bits_param : _GEN_40; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  assign io_out_bits_size = 3'h4 == chosen ? io_in_4_bits_size : _GEN_41; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  assign io_out_bits_source = 3'h4 == chosen ? io_in_4_bits_source : _GEN_42; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  assign io_out_bits_address = 3'h4 == chosen ? io_in_4_bits_address : 32'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  assign io_out_bits_data = 3'h4 == chosen ? io_in_4_bits_data : _GEN_44; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  assign io_out_bits_corrupt = 3'h4 == chosen ? io_in_4_bits_corrupt : _GEN_45; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  assign io_out_bits_union = 3'h4 == chosen ? io_in_4_bits_union : _GEN_46; // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  assign io_out_bits_last = 3'h4 == chosen ? io_in_4_bits_last : 3'h3 == chosen | (3'h2 == chosen | _GEN_23); // @[Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4 Arbiters.scala 42:16 chipyard.TestHarness.TinyRocketConfig.fir 185035:4]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiters.scala 25:20 chipyard.TestHarness.TinyRocketConfig.fir 185013:4]
      lockIdx <= 3'h0; // @[Arbiters.scala 25:20 chipyard.TestHarness.TinyRocketConfig.fir 185013:4]
    end else if (_T) begin // @[Arbiters.scala 58:24 chipyard.TestHarness.TinyRocketConfig.fir 185038:4]
      if (_T_1) begin // @[Arbiters.scala 59:50 chipyard.TestHarness.TinyRocketConfig.fir 185041:6]
        if (io_in_1_valid) begin // @[Mux.scala 47:69 chipyard.TestHarness.TinyRocketConfig.fir 185017:4]
          lockIdx <= 3'h1;
        end else begin
          lockIdx <= 3'h4;
        end
      end
    end
    if (reset) begin // @[Arbiters.scala 26:19 chipyard.TestHarness.TinyRocketConfig.fir 185014:4]
      locked <= 1'h0; // @[Arbiters.scala 26:19 chipyard.TestHarness.TinyRocketConfig.fir 185014:4]
    end else if (_T) begin // @[Arbiters.scala 58:24 chipyard.TestHarness.TinyRocketConfig.fir 185038:4]
      if (io_out_bits_last) begin // @[Arbiters.scala 64:35 chipyard.TestHarness.TinyRocketConfig.fir 185045:6]
        locked <= 1'h0; // @[Arbiters.scala 65:14 chipyard.TestHarness.TinyRocketConfig.fir 185046:8]
      end else begin
        locked <= _GEN_61;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockIdx = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  locked = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericSerializer_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 185050:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 185051:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 185052:4]
  output        io_in_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input         io_in_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input  [2:0]  io_in_bits_chanId, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input  [2:0]  io_in_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input  [2:0]  io_in_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input  [3:0]  io_in_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input  [1:0]  io_in_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input  [31:0] io_in_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input  [31:0] io_in_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input         io_in_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input  [3:0]  io_in_bits_union, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input         io_in_bits_last, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  input         io_out_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  output        io_out_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
  output [3:0]  io_out_bits // @[chipyard.TestHarness.TinyRocketConfig.fir 185053:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [84:0] data; // @[Serdes.scala 175:17 chipyard.TestHarness.TinyRocketConfig.fir 185055:4]
  reg  sending; // @[Serdes.scala 177:24 chipyard.TestHarness.TinyRocketConfig.fir 185056:4]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 185057:4]
  reg [4:0] sendCount; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 185058:4]
  wire  wrap_wrap = sendCount == 5'h15; // @[Counter.scala 72:24 chipyard.TestHarness.TinyRocketConfig.fir 185062:6]
  wire [4:0] _wrap_value_T_1 = sendCount + 5'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 185064:6]
  wire  sendDone = _T & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 185061:4 Counter.scala 118:24 chipyard.TestHarness.TinyRocketConfig.fir 185069:6 chipyard.TestHarness.TinyRocketConfig.fir 185060:4]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 185076:4]
  wire [84:0] _data_T = {io_in_bits_chanId,io_in_bits_opcode,io_in_bits_param,io_in_bits_size,io_in_bits_source,
    io_in_bits_address,io_in_bits_data,io_in_bits_corrupt,io_in_bits_union,io_in_bits_last}; // @[Serdes.scala 185:24 chipyard.TestHarness.TinyRocketConfig.fir 185086:6]
  wire  _GEN_4 = _T_1 | sending; // @[Serdes.scala 184:23 chipyard.TestHarness.TinyRocketConfig.fir 185077:4 Serdes.scala 186:13 chipyard.TestHarness.TinyRocketConfig.fir 185088:6 Serdes.scala 177:24 chipyard.TestHarness.TinyRocketConfig.fir 185056:4]
  wire [84:0] _data_T_1 = {{4'd0}, data[84:4]}; // @[Serdes.scala 189:39 chipyard.TestHarness.TinyRocketConfig.fir 185092:6]
  assign io_in_ready = ~sending; // @[Serdes.scala 180:18 chipyard.TestHarness.TinyRocketConfig.fir 185071:4]
  assign io_out_valid = sending; // @[Serdes.scala 181:16 chipyard.TestHarness.TinyRocketConfig.fir 185073:4]
  assign io_out_bits = data[3:0]; // @[Serdes.scala 182:22 chipyard.TestHarness.TinyRocketConfig.fir 185074:4]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 189:24 chipyard.TestHarness.TinyRocketConfig.fir 185091:4]
      data <= _data_T_1; // @[Serdes.scala 189:31 chipyard.TestHarness.TinyRocketConfig.fir 185093:6]
    end else if (_T_1) begin // @[Serdes.scala 184:23 chipyard.TestHarness.TinyRocketConfig.fir 185077:4]
      data <= _data_T; // @[Serdes.scala 185:10 chipyard.TestHarness.TinyRocketConfig.fir 185087:6]
    end
    if (reset) begin // @[Serdes.scala 177:24 chipyard.TestHarness.TinyRocketConfig.fir 185056:4]
      sending <= 1'h0; // @[Serdes.scala 177:24 chipyard.TestHarness.TinyRocketConfig.fir 185056:4]
    end else if (sendDone) begin // @[Serdes.scala 191:19 chipyard.TestHarness.TinyRocketConfig.fir 185095:4]
      sending <= 1'h0; // @[Serdes.scala 191:29 chipyard.TestHarness.TinyRocketConfig.fir 185096:6]
    end else begin
      sending <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 185058:4]
      sendCount <= 5'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 185058:4]
    end else if (_T) begin // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 185061:4]
      if (wrap_wrap) begin // @[Counter.scala 86:20 chipyard.TestHarness.TinyRocketConfig.fir 185066:6]
        sendCount <= 5'h0; // @[Counter.scala 86:28 chipyard.TestHarness.TinyRocketConfig.fir 185067:8]
      end else begin
        sendCount <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 185065:6]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  data = _RAND_0[84:0];
  _RAND_1 = {1{`RANDOM}};
  sending = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sendCount = _RAND_2[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericDeserializer_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 185099:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 185100:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 185101:4]
  output        io_in_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  input         io_in_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  input  [3:0]  io_in_bits, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  input         io_out_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  output        io_out_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  output [2:0]  io_out_bits_chanId, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  output [2:0]  io_out_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  output [2:0]  io_out_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  output [3:0]  io_out_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  output [1:0]  io_out_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  output [31:0] io_out_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  output [31:0] io_out_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  output        io_out_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
  output [3:0]  io_out_bits_union // @[chipyard.TestHarness.TinyRocketConfig.fir 185102:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] data_0; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_1; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_2; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_3; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_4; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_5; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_6; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_7; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_8; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_9; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_10; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_11; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_12; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_13; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_14; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_15; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_16; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_17; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_18; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_19; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_20; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg [3:0] data_21; // @[Serdes.scala 202:17 chipyard.TestHarness.TinyRocketConfig.fir 185104:4]
  reg  receiving; // @[Serdes.scala 204:26 chipyard.TestHarness.TinyRocketConfig.fir 185105:4]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 185106:4]
  reg [4:0] recvCount; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 185107:4]
  wire  wrap_wrap = recvCount == 5'h15; // @[Counter.scala 72:24 chipyard.TestHarness.TinyRocketConfig.fir 185111:6]
  wire [4:0] _wrap_value_T_1 = recvCount + 5'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 185113:6]
  wire  recvDone = _T & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 185110:4 Counter.scala 118:24 chipyard.TestHarness.TinyRocketConfig.fir 185118:6 chipyard.TestHarness.TinyRocketConfig.fir 185109:4]
  wire [19:0] io_out_bits_lo_lo = {data_4,data_3,data_2,data_1,data_0}; // @[Serdes.scala 209:23 chipyard.TestHarness.TinyRocketConfig.fir 185126:4]
  wire [43:0] io_out_bits_lo = {data_10,data_9,data_8,data_7,data_6,data_5,io_out_bits_lo_lo}; // @[Serdes.scala 209:23 chipyard.TestHarness.TinyRocketConfig.fir 185132:4]
  wire [19:0] io_out_bits_hi_lo = {data_15,data_14,data_13,data_12,data_11}; // @[Serdes.scala 209:23 chipyard.TestHarness.TinyRocketConfig.fir 185136:4]
  wire [87:0] _io_out_bits_T = {data_21,data_20,data_19,data_18,data_17,data_16,io_out_bits_hi_lo,io_out_bits_lo}; // @[Serdes.scala 209:23 chipyard.TestHarness.TinyRocketConfig.fir 185143:4]
  wire  _GEN_47 = recvDone ? 1'h0 : receiving; // @[Serdes.scala 215:19 chipyard.TestHarness.TinyRocketConfig.fir 185181:4 Serdes.scala 215:31 chipyard.TestHarness.TinyRocketConfig.fir 185182:6 Serdes.scala 204:26 chipyard.TestHarness.TinyRocketConfig.fir 185105:4]
  wire  _T_2 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 185184:4]
  wire  _GEN_48 = _T_2 | _GEN_47; // @[Serdes.scala 217:24 chipyard.TestHarness.TinyRocketConfig.fir 185185:4 Serdes.scala 217:36 chipyard.TestHarness.TinyRocketConfig.fir 185186:6]
  assign io_in_ready = receiving; // @[Serdes.scala 207:15 chipyard.TestHarness.TinyRocketConfig.fir 185120:4]
  assign io_out_valid = ~receiving; // @[Serdes.scala 208:19 chipyard.TestHarness.TinyRocketConfig.fir 185121:4]
  assign io_out_bits_chanId = _io_out_bits_T[84:82]; // @[Serdes.scala 209:38 chipyard.TestHarness.TinyRocketConfig.fir 185165:4]
  assign io_out_bits_opcode = _io_out_bits_T[81:79]; // @[Serdes.scala 209:38 chipyard.TestHarness.TinyRocketConfig.fir 185163:4]
  assign io_out_bits_param = _io_out_bits_T[78:76]; // @[Serdes.scala 209:38 chipyard.TestHarness.TinyRocketConfig.fir 185161:4]
  assign io_out_bits_size = _io_out_bits_T[75:72]; // @[Serdes.scala 209:38 chipyard.TestHarness.TinyRocketConfig.fir 185159:4]
  assign io_out_bits_source = _io_out_bits_T[71:70]; // @[Serdes.scala 209:38 chipyard.TestHarness.TinyRocketConfig.fir 185157:4]
  assign io_out_bits_address = _io_out_bits_T[69:38]; // @[Serdes.scala 209:38 chipyard.TestHarness.TinyRocketConfig.fir 185155:4]
  assign io_out_bits_data = _io_out_bits_T[37:6]; // @[Serdes.scala 209:38 chipyard.TestHarness.TinyRocketConfig.fir 185153:4]
  assign io_out_bits_corrupt = _io_out_bits_T[5]; // @[Serdes.scala 209:38 chipyard.TestHarness.TinyRocketConfig.fir 185151:4]
  assign io_out_bits_union = _io_out_bits_T[4:1]; // @[Serdes.scala 209:38 chipyard.TestHarness.TinyRocketConfig.fir 185149:4]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h0 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_0 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h1 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_1 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h2 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_2 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h3 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_3 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h4 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_4 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h5 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_5 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h6 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_6 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h7 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_7 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h8 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_8 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h9 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_9 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'ha == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_10 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'hb == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_11 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'hc == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_12 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'hd == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_13 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'he == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_14 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'hf == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_15 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h10 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_16 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h11 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_17 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h12 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_18 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h13 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_19 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h14 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_20 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.TinyRocketConfig.fir 185178:4]
      if (5'h15 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
        data_21 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 185179:6]
      end
    end
    receiving <= reset | _GEN_48; // @[Serdes.scala 204:26 chipyard.TestHarness.TinyRocketConfig.fir 185105:4 Serdes.scala 204:26 chipyard.TestHarness.TinyRocketConfig.fir 185105:4]
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 185107:4]
      recvCount <= 5'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 185107:4]
    end else if (_T) begin // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 185110:4]
      if (wrap_wrap) begin // @[Counter.scala 86:20 chipyard.TestHarness.TinyRocketConfig.fir 185115:6]
        recvCount <= 5'h0; // @[Counter.scala 86:28 chipyard.TestHarness.TinyRocketConfig.fir 185116:8]
      end else begin
        recvCount <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 185114:6]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  data_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  data_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  data_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  data_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  data_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  data_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  data_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  data_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  data_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  data_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  data_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  data_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  data_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  data_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  data_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  data_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  data_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  data_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  data_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  data_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  data_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  receiving = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  recvCount = _RAND_23[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SerialAdapter_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 195938:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 195939:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 195940:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 195941:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 195941:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 195941:4]
  output [3:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 195941:4]
  output [31:0] auto_out_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 195941:4]
  output [3:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 195941:4]
  output [31:0] auto_out_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 195941:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 195941:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 195941:4]
  input  [31:0] auto_out_d_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 195941:4]
  output        io_serial_in_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 195942:4]
  input         io_serial_in_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 195942:4]
  input  [31:0] io_serial_in_bits, // @[chipyard.TestHarness.TinyRocketConfig.fir 195942:4]
  input         io_serial_out_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 195942:4]
  output        io_serial_out_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 195942:4]
  output [31:0] io_serial_out_bits // @[chipyard.TestHarness.TinyRocketConfig.fir 195942:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cmd; // @[SerialAdapter.scala 86:16 chipyard.TestHarness.TinyRocketConfig.fir 195951:4]
  reg [63:0] addr; // @[SerialAdapter.scala 87:17 chipyard.TestHarness.TinyRocketConfig.fir 195952:4]
  reg [63:0] len; // @[SerialAdapter.scala 88:16 chipyard.TestHarness.TinyRocketConfig.fir 195953:4]
  reg [31:0] body_0; // @[SerialAdapter.scala 89:17 chipyard.TestHarness.TinyRocketConfig.fir 195954:4]
  reg  bodyValid; // @[SerialAdapter.scala 90:22 chipyard.TestHarness.TinyRocketConfig.fir 195955:4]
  reg  idx; // @[SerialAdapter.scala 91:16 chipyard.TestHarness.TinyRocketConfig.fir 195956:4]
  reg [3:0] state; // @[SerialAdapter.scala 97:22 chipyard.TestHarness.TinyRocketConfig.fir 195957:4]
  wire  _io_serial_in_ready_T = state == 4'h0; // @[package.scala 15:47 chipyard.TestHarness.TinyRocketConfig.fir 195958:4]
  wire  _io_serial_in_ready_T_1 = state == 4'h1; // @[package.scala 15:47 chipyard.TestHarness.TinyRocketConfig.fir 195959:4]
  wire  _io_serial_in_ready_T_2 = state == 4'h2; // @[package.scala 15:47 chipyard.TestHarness.TinyRocketConfig.fir 195960:4]
  wire  _io_serial_in_ready_T_3 = state == 4'h6; // @[package.scala 15:47 chipyard.TestHarness.TinyRocketConfig.fir 195961:4]
  wire  _io_serial_in_ready_T_4 = _io_serial_in_ready_T | _io_serial_in_ready_T_1; // @[package.scala 72:59 chipyard.TestHarness.TinyRocketConfig.fir 195962:4]
  wire  _io_serial_in_ready_T_5 = _io_serial_in_ready_T_4 | _io_serial_in_ready_T_2; // @[package.scala 72:59 chipyard.TestHarness.TinyRocketConfig.fir 195963:4]
  wire  _io_serial_out_valid_T = state == 4'h5; // @[SerialAdapter.scala 100:32 chipyard.TestHarness.TinyRocketConfig.fir 195966:4]
  wire [29:0] beatAddr = addr[31:2]; // @[SerialAdapter.scala 103:22 chipyard.TestHarness.TinyRocketConfig.fir 195969:4]
  wire [29:0] nextAddr_hi = beatAddr + 30'h1; // @[SerialAdapter.scala 104:31 chipyard.TestHarness.TinyRocketConfig.fir 195971:4]
  wire [31:0] nextAddr = {nextAddr_hi,2'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 195972:4]
  wire [3:0] wmask = bodyValid ? 4'hf : 4'h0; // @[Bitwise.scala 72:12 chipyard.TestHarness.TinyRocketConfig.fir 195975:4]
  wire [63:0] _GEN_49 = {{32'd0}, nextAddr}; // @[SerialAdapter.scala 107:28 chipyard.TestHarness.TinyRocketConfig.fir 195976:4]
  wire [63:0] addr_size = _GEN_49 - addr; // @[SerialAdapter.scala 107:28 chipyard.TestHarness.TinyRocketConfig.fir 195977:4]
  wire [63:0] len_size_hi = len + 64'h1; // @[SerialAdapter.scala 108:26 chipyard.TestHarness.TinyRocketConfig.fir 195979:4]
  wire [65:0] len_size = {len_size_hi,2'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 195980:4]
  wire [65:0] _GEN_50 = {{2'd0}, addr_size}; // @[SerialAdapter.scala 109:31 chipyard.TestHarness.TinyRocketConfig.fir 195981:4]
  wire  _raw_size_T = len_size < _GEN_50; // @[SerialAdapter.scala 109:31 chipyard.TestHarness.TinyRocketConfig.fir 195981:4]
  wire [65:0] raw_size = _raw_size_T ? len_size : {{2'd0}, addr_size}; // @[SerialAdapter.scala 109:21 chipyard.TestHarness.TinyRocketConfig.fir 195982:4]
  wire  _rsize_T = 66'h1 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.TinyRocketConfig.fir 195983:4]
  wire [1:0] _rsize_T_1 = _rsize_T ? 2'h0 : 2'h2; // @[Mux.scala 80:57 chipyard.TestHarness.TinyRocketConfig.fir 195984:4]
  wire  _rsize_T_2 = 66'h2 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.TinyRocketConfig.fir 195985:4]
  wire [1:0] rsize = _rsize_T_2 ? 2'h1 : _rsize_T_1; // @[Mux.scala 80:57 chipyard.TestHarness.TinyRocketConfig.fir 195986:4]
  wire [1:0] _pow2size_T_66 = raw_size[0] + raw_size[1]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196053:4]
  wire [1:0] _pow2size_T_68 = raw_size[2] + raw_size[3]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196055:4]
  wire [2:0] _pow2size_T_70 = _pow2size_T_66 + _pow2size_T_68; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196057:4]
  wire [1:0] _pow2size_T_72 = raw_size[4] + raw_size[5]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196059:4]
  wire [1:0] _pow2size_T_74 = raw_size[6] + raw_size[7]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196061:4]
  wire [2:0] _pow2size_T_76 = _pow2size_T_72 + _pow2size_T_74; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196063:4]
  wire [3:0] _pow2size_T_78 = _pow2size_T_70 + _pow2size_T_76; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196065:4]
  wire [1:0] _pow2size_T_80 = raw_size[8] + raw_size[9]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196067:4]
  wire [1:0] _pow2size_T_82 = raw_size[10] + raw_size[11]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196069:4]
  wire [2:0] _pow2size_T_84 = _pow2size_T_80 + _pow2size_T_82; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196071:4]
  wire [1:0] _pow2size_T_86 = raw_size[12] + raw_size[13]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196073:4]
  wire [1:0] _pow2size_T_88 = raw_size[14] + raw_size[15]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196075:4]
  wire [2:0] _pow2size_T_90 = _pow2size_T_86 + _pow2size_T_88; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196077:4]
  wire [3:0] _pow2size_T_92 = _pow2size_T_84 + _pow2size_T_90; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196079:4]
  wire [4:0] _pow2size_T_94 = _pow2size_T_78 + _pow2size_T_92; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196081:4]
  wire [1:0] _pow2size_T_96 = raw_size[16] + raw_size[17]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196083:4]
  wire [1:0] _pow2size_T_98 = raw_size[18] + raw_size[19]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196085:4]
  wire [2:0] _pow2size_T_100 = _pow2size_T_96 + _pow2size_T_98; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196087:4]
  wire [1:0] _pow2size_T_102 = raw_size[20] + raw_size[21]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196089:4]
  wire [1:0] _pow2size_T_104 = raw_size[22] + raw_size[23]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196091:4]
  wire [2:0] _pow2size_T_106 = _pow2size_T_102 + _pow2size_T_104; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196093:4]
  wire [3:0] _pow2size_T_108 = _pow2size_T_100 + _pow2size_T_106; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196095:4]
  wire [1:0] _pow2size_T_110 = raw_size[24] + raw_size[25]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196097:4]
  wire [1:0] _pow2size_T_112 = raw_size[26] + raw_size[27]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196099:4]
  wire [2:0] _pow2size_T_114 = _pow2size_T_110 + _pow2size_T_112; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196101:4]
  wire [1:0] _pow2size_T_116 = raw_size[28] + raw_size[29]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196103:4]
  wire [1:0] _pow2size_T_118 = raw_size[31] + raw_size[32]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196105:4]
  wire [1:0] _GEN_51 = {{1'd0}, raw_size[30]}; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196107:4]
  wire [2:0] _pow2size_T_120 = _GEN_51 + _pow2size_T_118; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196107:4]
  wire [2:0] _pow2size_T_122 = _pow2size_T_116 + _pow2size_T_120[1:0]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196109:4]
  wire [3:0] _pow2size_T_124 = _pow2size_T_114 + _pow2size_T_122; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196111:4]
  wire [4:0] _pow2size_T_126 = _pow2size_T_108 + _pow2size_T_124; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196113:4]
  wire [5:0] _pow2size_T_128 = _pow2size_T_94 + _pow2size_T_126; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196115:4]
  wire [1:0] _pow2size_T_130 = raw_size[33] + raw_size[34]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196117:4]
  wire [1:0] _pow2size_T_132 = raw_size[35] + raw_size[36]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196119:4]
  wire [2:0] _pow2size_T_134 = _pow2size_T_130 + _pow2size_T_132; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196121:4]
  wire [1:0] _pow2size_T_136 = raw_size[37] + raw_size[38]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196123:4]
  wire [1:0] _pow2size_T_138 = raw_size[39] + raw_size[40]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196125:4]
  wire [2:0] _pow2size_T_140 = _pow2size_T_136 + _pow2size_T_138; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196127:4]
  wire [3:0] _pow2size_T_142 = _pow2size_T_134 + _pow2size_T_140; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196129:4]
  wire [1:0] _pow2size_T_144 = raw_size[41] + raw_size[42]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196131:4]
  wire [1:0] _pow2size_T_146 = raw_size[43] + raw_size[44]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196133:4]
  wire [2:0] _pow2size_T_148 = _pow2size_T_144 + _pow2size_T_146; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196135:4]
  wire [1:0] _pow2size_T_150 = raw_size[45] + raw_size[46]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196137:4]
  wire [1:0] _pow2size_T_152 = raw_size[47] + raw_size[48]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196139:4]
  wire [2:0] _pow2size_T_154 = _pow2size_T_150 + _pow2size_T_152; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196141:4]
  wire [3:0] _pow2size_T_156 = _pow2size_T_148 + _pow2size_T_154; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196143:4]
  wire [4:0] _pow2size_T_158 = _pow2size_T_142 + _pow2size_T_156; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196145:4]
  wire [1:0] _pow2size_T_160 = raw_size[49] + raw_size[50]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196147:4]
  wire [1:0] _pow2size_T_162 = raw_size[51] + raw_size[52]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196149:4]
  wire [2:0] _pow2size_T_164 = _pow2size_T_160 + _pow2size_T_162; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196151:4]
  wire [1:0] _pow2size_T_166 = raw_size[53] + raw_size[54]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196153:4]
  wire [1:0] _pow2size_T_168 = raw_size[55] + raw_size[56]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196155:4]
  wire [2:0] _pow2size_T_170 = _pow2size_T_166 + _pow2size_T_168; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196157:4]
  wire [3:0] _pow2size_T_172 = _pow2size_T_164 + _pow2size_T_170; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196159:4]
  wire [1:0] _pow2size_T_174 = raw_size[57] + raw_size[58]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196161:4]
  wire [1:0] _pow2size_T_176 = raw_size[59] + raw_size[60]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196163:4]
  wire [2:0] _pow2size_T_178 = _pow2size_T_174 + _pow2size_T_176; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196165:4]
  wire [1:0] _pow2size_T_180 = raw_size[61] + raw_size[62]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196167:4]
  wire [1:0] _pow2size_T_182 = raw_size[64] + raw_size[65]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196169:4]
  wire [1:0] _GEN_52 = {{1'd0}, raw_size[63]}; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196171:4]
  wire [2:0] _pow2size_T_184 = _GEN_52 + _pow2size_T_182; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196171:4]
  wire [2:0] _pow2size_T_186 = _pow2size_T_180 + _pow2size_T_184[1:0]; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196173:4]
  wire [3:0] _pow2size_T_188 = _pow2size_T_178 + _pow2size_T_186; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196175:4]
  wire [4:0] _pow2size_T_190 = _pow2size_T_172 + _pow2size_T_188; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196177:4]
  wire [5:0] _pow2size_T_192 = _pow2size_T_158 + _pow2size_T_190; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196179:4]
  wire [6:0] _pow2size_T_194 = _pow2size_T_128 + _pow2size_T_192; // @[Bitwise.scala 47:55 chipyard.TestHarness.TinyRocketConfig.fir 196181:4]
  wire  pow2size = _pow2size_T_194 == 7'h1; // @[SerialAdapter.scala 113:37 chipyard.TestHarness.TinyRocketConfig.fir 196183:4]
  wire [1:0] byteAddr = pow2size ? addr[1:0] : 2'h0; // @[SerialAdapter.scala 114:21 chipyard.TestHarness.TinyRocketConfig.fir 196185:4]
  wire [31:0] _GEN_53 = {beatAddr, 2'h0}; // @[SerialAdapter.scala 117:19 chipyard.TestHarness.TinyRocketConfig.fir 196186:4]
  wire [32:0] _put_acquire_T = {{1'd0}, _GEN_53}; // @[SerialAdapter.scala 117:19 chipyard.TestHarness.TinyRocketConfig.fir 196186:4]
  wire [31:0] get_acquire_address = {beatAddr,byteAddr}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 196251:4]
  wire  get_acquire_a_mask_sizeOH_shiftAmount = rsize[0]; // @[OneHot.scala 64:49 chipyard.TestHarness.TinyRocketConfig.fir 196312:4]
  wire [1:0] _get_acquire_a_mask_sizeOH_T_1 = 2'h1 << get_acquire_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.TinyRocketConfig.fir 196313:4]
  wire [1:0] get_acquire_a_mask_sizeOH = _get_acquire_a_mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81 chipyard.TestHarness.TinyRocketConfig.fir 196315:4]
  wire  _get_acquire_a_mask_T = rsize >= 2'h2; // @[Misc.scala 205:21 chipyard.TestHarness.TinyRocketConfig.fir 196316:4]
  wire  get_acquire_a_mask_size = get_acquire_a_mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 196317:4]
  wire  get_acquire_a_mask_bit = get_acquire_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 196318:4]
  wire  get_acquire_a_mask_nbit = ~get_acquire_a_mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 196319:4]
  wire  _get_acquire_a_mask_acc_T = get_acquire_a_mask_size & get_acquire_a_mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196321:4]
  wire  get_acquire_a_mask_acc = _get_acquire_a_mask_T | _get_acquire_a_mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196322:4]
  wire  _get_acquire_a_mask_acc_T_1 = get_acquire_a_mask_size & get_acquire_a_mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196324:4]
  wire  get_acquire_a_mask_acc_1 = _get_acquire_a_mask_T | _get_acquire_a_mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196325:4]
  wire  get_acquire_a_mask_size_1 = get_acquire_a_mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 196326:4]
  wire  get_acquire_a_mask_bit_1 = get_acquire_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 196327:4]
  wire  get_acquire_a_mask_nbit_1 = ~get_acquire_a_mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 196328:4]
  wire  get_acquire_a_mask_eq_2 = get_acquire_a_mask_nbit & get_acquire_a_mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 196329:4]
  wire  _get_acquire_a_mask_acc_T_2 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196330:4]
  wire  get_acquire_a_mask_lo_lo = get_acquire_a_mask_acc | _get_acquire_a_mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196331:4]
  wire  get_acquire_a_mask_eq_3 = get_acquire_a_mask_nbit & get_acquire_a_mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 196332:4]
  wire  _get_acquire_a_mask_acc_T_3 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196333:4]
  wire  get_acquire_a_mask_lo_hi = get_acquire_a_mask_acc | _get_acquire_a_mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196334:4]
  wire  get_acquire_a_mask_eq_4 = get_acquire_a_mask_bit & get_acquire_a_mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 196335:4]
  wire  _get_acquire_a_mask_acc_T_4 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196336:4]
  wire  get_acquire_a_mask_hi_lo = get_acquire_a_mask_acc_1 | _get_acquire_a_mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196337:4]
  wire  get_acquire_a_mask_eq_5 = get_acquire_a_mask_bit & get_acquire_a_mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 196338:4]
  wire  _get_acquire_a_mask_acc_T_5 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196339:4]
  wire  get_acquire_a_mask_hi_hi = get_acquire_a_mask_acc_1 | _get_acquire_a_mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196340:4]
  wire [3:0] get_acquire_mask = {get_acquire_a_mask_hi_hi,get_acquire_a_mask_hi_lo,get_acquire_a_mask_lo_hi,
    get_acquire_a_mask_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 196343:4]
  wire  _bundleOut_0_a_valid_T = state == 4'h7; // @[package.scala 15:47 chipyard.TestHarness.TinyRocketConfig.fir 196347:4]
  wire  _bundleOut_0_a_valid_T_1 = state == 4'h3; // @[package.scala 15:47 chipyard.TestHarness.TinyRocketConfig.fir 196348:4]
  wire [3:0] get_acquire_size = {{2'd0}, rsize}; // @[Edges.scala 447:17 chipyard.TestHarness.TinyRocketConfig.fir 196304:4 Edges.scala 450:15 chipyard.TestHarness.TinyRocketConfig.fir 196308:4]
  wire [31:0] put_acquire_address = _put_acquire_T[31:0]; // @[Edges.scala 483:17 chipyard.TestHarness.TinyRocketConfig.fir 196241:4 Edges.scala 488:15 chipyard.TestHarness.TinyRocketConfig.fir 196247:4]
  wire  _bundleOut_0_d_ready_T = state == 4'h8; // @[package.scala 15:47 chipyard.TestHarness.TinyRocketConfig.fir 196367:4]
  wire  _bundleOut_0_d_ready_T_1 = state == 4'h4; // @[package.scala 15:47 chipyard.TestHarness.TinyRocketConfig.fir 196368:4]
  wire  _T_1 = _io_serial_in_ready_T & io_serial_in_valid; // @[SerialAdapter.scala 138:25 chipyard.TestHarness.TinyRocketConfig.fir 196375:4]
  wire  _GEN_1 = _T_1 ? 1'h0 : idx; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.TinyRocketConfig.fir 196376:4 SerialAdapter.scala 140:9 chipyard.TestHarness.TinyRocketConfig.fir 196378:6 SerialAdapter.scala 91:16 chipyard.TestHarness.TinyRocketConfig.fir 195956:4]
  wire [63:0] _GEN_2 = _T_1 ? 64'h0 : addr; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.TinyRocketConfig.fir 196376:4 SerialAdapter.scala 141:10 chipyard.TestHarness.TinyRocketConfig.fir 196379:6 SerialAdapter.scala 87:17 chipyard.TestHarness.TinyRocketConfig.fir 195952:4]
  wire [63:0] _GEN_3 = _T_1 ? 64'h0 : len; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.TinyRocketConfig.fir 196376:4 SerialAdapter.scala 142:9 chipyard.TestHarness.TinyRocketConfig.fir 196380:6 SerialAdapter.scala 88:16 chipyard.TestHarness.TinyRocketConfig.fir 195953:4]
  wire [3:0] _GEN_4 = _T_1 ? 4'h1 : state; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.TinyRocketConfig.fir 196376:4 SerialAdapter.scala 143:11 chipyard.TestHarness.TinyRocketConfig.fir 196381:6 SerialAdapter.scala 97:22 chipyard.TestHarness.TinyRocketConfig.fir 195957:4]
  wire  _T_3 = _io_serial_in_ready_T_1 & io_serial_in_valid; // @[SerialAdapter.scala 146:26 chipyard.TestHarness.TinyRocketConfig.fir 196384:4]
  wire [5:0] _addr_T = {idx,5'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 196387:6]
  wire [94:0] _GEN_54 = {{63'd0}, io_serial_in_bits}; // @[SerialAdapter.scala 132:12 chipyard.TestHarness.TinyRocketConfig.fir 196388:6]
  wire [94:0] _addr_T_1 = _GEN_54 << _addr_T; // @[SerialAdapter.scala 132:12 chipyard.TestHarness.TinyRocketConfig.fir 196388:6]
  wire [94:0] _GEN_55 = {{31'd0}, addr}; // @[SerialAdapter.scala 147:18 chipyard.TestHarness.TinyRocketConfig.fir 196389:6]
  wire [94:0] _addr_T_2 = _GEN_55 | _addr_T_1; // @[SerialAdapter.scala 147:18 chipyard.TestHarness.TinyRocketConfig.fir 196389:6]
  wire  _idx_T_1 = idx + 1'h1; // @[SerialAdapter.scala 148:16 chipyard.TestHarness.TinyRocketConfig.fir 196392:6]
  wire  _GEN_5 = idx ? 1'h0 : _idx_T_1; // @[SerialAdapter.scala 149:43 chipyard.TestHarness.TinyRocketConfig.fir 196395:6 SerialAdapter.scala 150:11 chipyard.TestHarness.TinyRocketConfig.fir 196396:8 SerialAdapter.scala 148:9 chipyard.TestHarness.TinyRocketConfig.fir 196393:6]
  wire [3:0] _GEN_6 = idx ? 4'h2 : _GEN_4; // @[SerialAdapter.scala 149:43 chipyard.TestHarness.TinyRocketConfig.fir 196395:6 SerialAdapter.scala 151:13 chipyard.TestHarness.TinyRocketConfig.fir 196397:8]
  wire [94:0] _GEN_7 = _T_3 ? _addr_T_2 : {{31'd0}, _GEN_2}; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.TinyRocketConfig.fir 196385:4 SerialAdapter.scala 147:10 chipyard.TestHarness.TinyRocketConfig.fir 196390:6]
  wire  _GEN_8 = _T_3 ? _GEN_5 : _GEN_1; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.TinyRocketConfig.fir 196385:4]
  wire [3:0] _GEN_9 = _T_3 ? _GEN_6 : _GEN_4; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.TinyRocketConfig.fir 196385:4]
  wire  _T_6 = _io_serial_in_ready_T_2 & io_serial_in_valid; // @[SerialAdapter.scala 155:25 chipyard.TestHarness.TinyRocketConfig.fir 196401:4]
  wire [94:0] _GEN_57 = {{31'd0}, len}; // @[SerialAdapter.scala 156:16 chipyard.TestHarness.TinyRocketConfig.fir 196406:6]
  wire [94:0] _len_T_2 = _GEN_57 | _addr_T_1; // @[SerialAdapter.scala 156:16 chipyard.TestHarness.TinyRocketConfig.fir 196406:6]
  wire  _T_8 = cmd == 32'h1; // @[SerialAdapter.scala 160:17 chipyard.TestHarness.TinyRocketConfig.fir 196414:8]
  wire  _T_9 = cmd == 32'h0; // @[SerialAdapter.scala 163:24 chipyard.TestHarness.TinyRocketConfig.fir 196420:10]
  wire  _T_12 = ~reset; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.TinyRocketConfig.fir 196427:12]
  wire [3:0] _GEN_10 = _T_9 ? 4'h3 : _GEN_9; // @[SerialAdapter.scala 163:38 chipyard.TestHarness.TinyRocketConfig.fir 196421:10 SerialAdapter.scala 164:15 chipyard.TestHarness.TinyRocketConfig.fir 196422:12]
  wire  _GEN_11 = _T_8 ? 1'h0 : bodyValid; // @[SerialAdapter.scala 160:32 chipyard.TestHarness.TinyRocketConfig.fir 196415:8 SerialAdapter.scala 161:19 chipyard.TestHarness.TinyRocketConfig.fir 196416:10 SerialAdapter.scala 90:22 chipyard.TestHarness.TinyRocketConfig.fir 195955:4]
  wire [3:0] _GEN_12 = _T_8 ? 4'h6 : _GEN_10; // @[SerialAdapter.scala 160:32 chipyard.TestHarness.TinyRocketConfig.fir 196415:8 SerialAdapter.scala 162:15 chipyard.TestHarness.TinyRocketConfig.fir 196417:10]
  wire  _GEN_14 = idx ? _GEN_11 : bodyValid; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.TinyRocketConfig.fir 196412:6 SerialAdapter.scala 90:22 chipyard.TestHarness.TinyRocketConfig.fir 195955:4]
  wire [3:0] _GEN_15 = idx ? _GEN_12 : _GEN_9; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.TinyRocketConfig.fir 196412:6]
  wire [94:0] _GEN_16 = _T_6 ? _len_T_2 : {{31'd0}, _GEN_3}; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.TinyRocketConfig.fir 196402:4 SerialAdapter.scala 156:9 chipyard.TestHarness.TinyRocketConfig.fir 196407:6]
  wire  _GEN_17 = _T_6 ? _GEN_5 : _GEN_8; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.TinyRocketConfig.fir 196402:4]
  wire  _GEN_18 = _T_6 ? _GEN_14 : bodyValid; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.TinyRocketConfig.fir 196402:4 SerialAdapter.scala 90:22 chipyard.TestHarness.TinyRocketConfig.fir 195955:4]
  wire [3:0] _GEN_19 = _T_6 ? _GEN_15 : _GEN_9; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.TinyRocketConfig.fir 196402:4]
  wire  _T_14 = _bundleOut_0_a_valid_T_1 & auto_out_a_ready; // @[SerialAdapter.scala 171:30 chipyard.TestHarness.TinyRocketConfig.fir 196436:4]
  wire [3:0] _GEN_20 = _T_14 ? 4'h4 : _GEN_19; // @[SerialAdapter.scala 171:46 chipyard.TestHarness.TinyRocketConfig.fir 196437:4 SerialAdapter.scala 172:11 chipyard.TestHarness.TinyRocketConfig.fir 196438:6]
  wire  _T_16 = _bundleOut_0_d_ready_T_1 & auto_out_d_valid; // @[SerialAdapter.scala 175:31 chipyard.TestHarness.TinyRocketConfig.fir 196441:4]
  wire  _GEN_22 = _T_16 ? 1'h0 : _GEN_17; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.TinyRocketConfig.fir 196442:4 SerialAdapter.scala 177:9 chipyard.TestHarness.TinyRocketConfig.fir 196449:6]
  wire [94:0] _GEN_23 = _T_16 ? {{63'd0}, nextAddr} : _GEN_7; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.TinyRocketConfig.fir 196442:4 SerialAdapter.scala 178:10 chipyard.TestHarness.TinyRocketConfig.fir 196450:6]
  wire [3:0] _GEN_24 = _T_16 ? 4'h5 : _GEN_20; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.TinyRocketConfig.fir 196442:4 SerialAdapter.scala 179:11 chipyard.TestHarness.TinyRocketConfig.fir 196451:6]
  wire  _T_19 = _io_serial_out_valid_T & io_serial_out_ready; // @[SerialAdapter.scala 182:31 chipyard.TestHarness.TinyRocketConfig.fir 196454:4]
  wire [63:0] _len_T_4 = len - 64'h1; // @[SerialAdapter.scala 184:16 chipyard.TestHarness.TinyRocketConfig.fir 196460:6]
  wire  _T_20 = len == 64'h0; // @[SerialAdapter.scala 185:15 chipyard.TestHarness.TinyRocketConfig.fir 196462:6]
  wire  _T_21 = ~idx; // @[SerialAdapter.scala 186:20 chipyard.TestHarness.TinyRocketConfig.fir 196467:8]
  wire [3:0] _GEN_25 = _T_21 ? 4'h3 : _GEN_24; // @[SerialAdapter.scala 186:48 chipyard.TestHarness.TinyRocketConfig.fir 196468:8 SerialAdapter.scala 186:56 chipyard.TestHarness.TinyRocketConfig.fir 196469:10]
  wire [3:0] _GEN_26 = _T_20 ? 4'h0 : _GEN_25; // @[SerialAdapter.scala 185:24 chipyard.TestHarness.TinyRocketConfig.fir 196463:6 SerialAdapter.scala 185:32 chipyard.TestHarness.TinyRocketConfig.fir 196464:8]
  wire  _GEN_27 = _T_19 ? _idx_T_1 : _GEN_22; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.TinyRocketConfig.fir 196455:4 SerialAdapter.scala 183:9 chipyard.TestHarness.TinyRocketConfig.fir 196458:6]
  wire [94:0] _GEN_28 = _T_19 ? {{31'd0}, _len_T_4} : _GEN_16; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.TinyRocketConfig.fir 196455:4 SerialAdapter.scala 184:9 chipyard.TestHarness.TinyRocketConfig.fir 196461:6]
  wire [3:0] _GEN_29 = _T_19 ? _GEN_26 : _GEN_24; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.TinyRocketConfig.fir 196455:4]
  wire  _T_23 = _io_serial_in_ready_T_3 & io_serial_in_valid; // @[SerialAdapter.scala 189:32 chipyard.TestHarness.TinyRocketConfig.fir 196473:4]
  wire [1:0] _bodyValid_T = 2'h1 << idx; // @[OneHot.scala 58:35 chipyard.TestHarness.TinyRocketConfig.fir 196476:6]
  wire [1:0] _GEN_58 = {{1'd0}, bodyValid}; // @[SerialAdapter.scala 191:28 chipyard.TestHarness.TinyRocketConfig.fir 196477:6]
  wire [1:0] _bodyValid_T_1 = _GEN_58 | _bodyValid_T; // @[SerialAdapter.scala 191:28 chipyard.TestHarness.TinyRocketConfig.fir 196477:6]
  wire  _T_26 = _T_21 | _T_20; // @[SerialAdapter.scala 192:42 chipyard.TestHarness.TinyRocketConfig.fir 196481:6]
  wire [3:0] _GEN_30 = _T_26 ? 4'h7 : _GEN_29; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.TinyRocketConfig.fir 196482:6 SerialAdapter.scala 193:13 chipyard.TestHarness.TinyRocketConfig.fir 196483:8]
  wire  _GEN_31 = _T_26 ? _GEN_27 : _idx_T_1; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.TinyRocketConfig.fir 196482:6 SerialAdapter.scala 195:11 chipyard.TestHarness.TinyRocketConfig.fir 196488:8]
  wire [94:0] _GEN_32 = _T_26 ? _GEN_28 : {{31'd0}, _len_T_4}; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.TinyRocketConfig.fir 196482:6 SerialAdapter.scala 196:11 chipyard.TestHarness.TinyRocketConfig.fir 196491:8]
  wire [1:0] _GEN_34 = _T_23 ? _bodyValid_T_1 : {{1'd0}, _GEN_18}; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.TinyRocketConfig.fir 196474:4 SerialAdapter.scala 191:15 chipyard.TestHarness.TinyRocketConfig.fir 196478:6]
  wire  _GEN_36 = _T_23 ? _GEN_31 : _GEN_27; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.TinyRocketConfig.fir 196474:4]
  wire [94:0] _GEN_37 = _T_23 ? _GEN_32 : _GEN_28; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.TinyRocketConfig.fir 196474:4]
  wire  _T_28 = _bundleOut_0_a_valid_T & auto_out_a_ready; // @[SerialAdapter.scala 200:32 chipyard.TestHarness.TinyRocketConfig.fir 196495:4]
  wire  _T_30 = _bundleOut_0_d_ready_T & auto_out_d_valid; // @[SerialAdapter.scala 204:31 chipyard.TestHarness.TinyRocketConfig.fir 196500:4]
  wire [94:0] _GEN_40 = _T_20 ? _GEN_23 : {{63'd0}, nextAddr}; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.TinyRocketConfig.fir 196503:6 SerialAdapter.scala 208:12 chipyard.TestHarness.TinyRocketConfig.fir 196507:8]
  wire [94:0] _GEN_41 = _T_20 ? _GEN_37 : {{31'd0}, _len_T_4}; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.TinyRocketConfig.fir 196503:6 SerialAdapter.scala 209:11 chipyard.TestHarness.TinyRocketConfig.fir 196510:8]
  wire  _GEN_42 = _T_20 & _GEN_36; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.TinyRocketConfig.fir 196503:6 SerialAdapter.scala 210:11 chipyard.TestHarness.TinyRocketConfig.fir 196511:8]
  wire [1:0] _GEN_43 = _T_20 ? _GEN_34 : 2'h0; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.TinyRocketConfig.fir 196503:6 SerialAdapter.scala 211:17 chipyard.TestHarness.TinyRocketConfig.fir 196512:8]
  wire [94:0] _GEN_45 = _T_30 ? _GEN_40 : _GEN_23; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.TinyRocketConfig.fir 196501:4]
  wire [94:0] _GEN_46 = _T_30 ? _GEN_41 : _GEN_37; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.TinyRocketConfig.fir 196501:4]
  wire [1:0] _GEN_48 = _T_30 ? _GEN_43 : _GEN_34; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.TinyRocketConfig.fir 196501:4]
  wire  _GEN_63 = _T_6 & idx & ~_T_8 & ~_T_9; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.TinyRocketConfig.fir 196429:14]
  assign auto_out_a_valid = _bundleOut_0_a_valid_T | _bundleOut_0_a_valid_T_1; // @[package.scala 72:59 chipyard.TestHarness.TinyRocketConfig.fir 196349:4]
  assign auto_out_a_bits_opcode = _bundleOut_0_a_valid_T ? 3'h1 : 3'h4; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.TinyRocketConfig.fir 196352:4]
  assign auto_out_a_bits_size = _bundleOut_0_a_valid_T ? 4'h2 : get_acquire_size; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.TinyRocketConfig.fir 196352:4]
  assign auto_out_a_bits_address = _bundleOut_0_a_valid_T ? put_acquire_address : get_acquire_address; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.TinyRocketConfig.fir 196352:4]
  assign auto_out_a_bits_mask = _bundleOut_0_a_valid_T ? wmask : get_acquire_mask; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.TinyRocketConfig.fir 196352:4]
  assign auto_out_a_bits_data = _bundleOut_0_a_valid_T ? body_0 : 32'h0; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.TinyRocketConfig.fir 196352:4]
  assign auto_out_d_ready = _bundleOut_0_d_ready_T | _bundleOut_0_d_ready_T_1; // @[package.scala 72:59 chipyard.TestHarness.TinyRocketConfig.fir 196369:4]
  assign io_serial_in_ready = _io_serial_in_ready_T_5 | _io_serial_in_ready_T_3; // @[package.scala 72:59 chipyard.TestHarness.TinyRocketConfig.fir 195964:4]
  assign io_serial_out_valid = state == 4'h5; // @[SerialAdapter.scala 100:32 chipyard.TestHarness.TinyRocketConfig.fir 195966:4]
  assign io_serial_out_bits = body_0; // @[SerialAdapter.scala 101:22 chipyard.TestHarness.TinyRocketConfig.fir 195968:4]
  always @(posedge clock) begin
    if (_T_1) begin // @[SerialAdapter.scala 138:48 chipyard.TestHarness.TinyRocketConfig.fir 196376:4]
      cmd <= io_serial_in_bits; // @[SerialAdapter.scala 139:9 chipyard.TestHarness.TinyRocketConfig.fir 196377:6]
    end
    addr <= _GEN_45[63:0];
    len <= _GEN_46[63:0];
    if (_T_23) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.TinyRocketConfig.fir 196474:4]
      body_0 <= io_serial_in_bits; // @[SerialAdapter.scala 190:15 chipyard.TestHarness.TinyRocketConfig.fir 196475:6]
    end else if (_T_16) begin // @[SerialAdapter.scala 175:47 chipyard.TestHarness.TinyRocketConfig.fir 196442:4]
      body_0 <= auto_out_d_bits_data; // @[SerialAdapter.scala 176:10 chipyard.TestHarness.TinyRocketConfig.fir 196448:6]
    end
    bodyValid <= _GEN_48[0];
    if (_T_30) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.TinyRocketConfig.fir 196501:4]
      idx <= _GEN_42;
    end else if (_T_23) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.TinyRocketConfig.fir 196474:4]
      if (_T_26) begin // @[SerialAdapter.scala 192:58 chipyard.TestHarness.TinyRocketConfig.fir 196482:6]
        idx <= _GEN_27;
      end else begin
        idx <= _idx_T_1; // @[SerialAdapter.scala 195:11 chipyard.TestHarness.TinyRocketConfig.fir 196488:8]
      end
    end else begin
      idx <= _GEN_27;
    end
    if (reset) begin // @[SerialAdapter.scala 97:22 chipyard.TestHarness.TinyRocketConfig.fir 195957:4]
      state <= 4'h0; // @[SerialAdapter.scala 97:22 chipyard.TestHarness.TinyRocketConfig.fir 195957:4]
    end else if (_T_30) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.TinyRocketConfig.fir 196501:4]
      if (_T_20) begin // @[SerialAdapter.scala 205:24 chipyard.TestHarness.TinyRocketConfig.fir 196503:6]
        state <= 4'h0; // @[SerialAdapter.scala 206:13 chipyard.TestHarness.TinyRocketConfig.fir 196504:8]
      end else begin
        state <= 4'h6; // @[SerialAdapter.scala 212:13 chipyard.TestHarness.TinyRocketConfig.fir 196513:8]
      end
    end else if (_T_28) begin // @[SerialAdapter.scala 200:48 chipyard.TestHarness.TinyRocketConfig.fir 196496:4]
      state <= 4'h8; // @[SerialAdapter.scala 201:11 chipyard.TestHarness.TinyRocketConfig.fir 196497:6]
    end else if (_T_23) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.TinyRocketConfig.fir 196474:4]
      state <= _GEN_30;
    end else begin
      state <= _GEN_29;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & idx & ~_T_8 & ~_T_9 & _T_12) begin
          $fwrite(32'h80000002,
            "Assertion failed: Bad TSI command\n    at SerialAdapter.scala:166 assert(false.B, \"Bad TSI command\")\n"); // @[SerialAdapter.scala 166:15 chipyard.TestHarness.TinyRocketConfig.fir 196429:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_63 & _T_12) begin
          $fatal; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.TinyRocketConfig.fir 196430:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cmd = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  addr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  len = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  body_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  bodyValid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  idx = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_41_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 196533:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 196534:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 196535:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input  [3:0]  io_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input         io_in_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input  [31:0] io_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input  [3:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input  [3:0]  io_in_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input         io_in_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input         io_in_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 196536:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 198373:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 198680:4]
  wire  _source_ok_T = ~io_in_a_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.TinyRocketConfig.fir 196547:6]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 196552:6]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 196554:6]
  wire [31:0] _GEN_71 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.TinyRocketConfig.fir 196555:6]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.TinyRocketConfig.fir 196555:6]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24 chipyard.TestHarness.TinyRocketConfig.fir 196556:6]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49 chipyard.TestHarness.TinyRocketConfig.fir 196558:6]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.TinyRocketConfig.fir 196559:6]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81 chipyard.TestHarness.TinyRocketConfig.fir 196561:6]
  wire  _mask_T = io_in_a_bits_size >= 4'h2; // @[Misc.scala 205:21 chipyard.TestHarness.TinyRocketConfig.fir 196562:6]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 196563:6]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 196564:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 196565:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196567:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196568:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196570:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196571:6]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 196572:6]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 196573:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 196574:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 196575:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196576:6]
  wire  mask_lo_lo = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196577:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 196578:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196579:6]
  wire  mask_lo_hi = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196580:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 196581:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196582:6]
  wire  mask_hi_lo = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196583:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 196584:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 196585:6]
  wire  mask_hi_hi = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 196586:6]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 196589:6]
  wire [32:0] _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 196593:6]
  wire  _T_15 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.TinyRocketConfig.fir 196605:6]
  wire  _T_17 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42 chipyard.TestHarness.TinyRocketConfig.fir 196608:8]
  wire  _T_20 = _T_17 & _source_ok_T; // @[Parameters.scala 1160:30 chipyard.TestHarness.TinyRocketConfig.fir 196611:8]
  wire [32:0] _T_26 = $signed(_T_7) & -33'sh101000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 196617:8]
  wire  _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 196618:8]
  wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 196619:8]
  wire [32:0] _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 196620:8]
  wire [32:0] _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 196622:8]
  wire  _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 196623:8]
  wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 196624:8]
  wire [32:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 196625:8]
  wire [32:0] _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 196627:8]
  wire  _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 196628:8]
  wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 196629:8]
  wire [32:0] _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 196630:8]
  wire [32:0] _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 196632:8]
  wire  _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 196633:8]
  wire [31:0] _T_43 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 196634:8]
  wire [32:0] _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 196635:8]
  wire [32:0] _T_46 = $signed(_T_44) & -33'sh4000000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 196637:8]
  wire  _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 196638:8]
  wire [31:0] _T_48 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 196639:8]
  wire [32:0] _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 196640:8]
  wire [32:0] _T_51 = $signed(_T_49) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 196642:8]
  wire  _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 196643:8]
  wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h54000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 196644:8]
  wire [32:0] _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 196645:8]
  wire [32:0] _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 196647:8]
  wire  _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 196648:8]
  wire [31:0] _T_58 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 196649:8]
  wire [32:0] _T_59 = {1'b0,$signed(_T_58)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 196650:8]
  wire [32:0] _T_61 = $signed(_T_59) & -33'sh4000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 196652:8]
  wire  _T_62 = $signed(_T_61) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 196653:8]
  wire  _T_63 = _T_27 | _T_32; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 196654:8]
  wire  _T_75 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196666:8]
  wire  _T_134 = _source_ok_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196733:8]
  wire  _T_135 = ~_T_134; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196734:8]
  wire  _T_138 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196741:8]
  wire  _T_139 = ~_T_138; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196742:8]
  wire  _T_141 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196748:8]
  wire  _T_142 = ~_T_141; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196749:8]
  wire  _T_143 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.TinyRocketConfig.fir 196754:8]
  wire  _T_145 = _T_143 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196756:8]
  wire  _T_146 = ~_T_145; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196757:8]
  wire [3:0] _T_147 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.TinyRocketConfig.fir 196762:8]
  wire  _T_148 = _T_147 == 4'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.TinyRocketConfig.fir 196763:8]
  wire  _T_150 = _T_148 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196765:8]
  wire  _T_151 = ~_T_150; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196766:8]
  wire  _T_152 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.TinyRocketConfig.fir 196771:8]
  wire  _T_154 = _T_152 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196773:8]
  wire  _T_155 = ~_T_154; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196774:8]
  wire  _T_156 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.TinyRocketConfig.fir 196780:6]
  wire  _T_288 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.TinyRocketConfig.fir 196937:8]
  wire  _T_290 = _T_288 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196939:8]
  wire  _T_291 = ~_T_290; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196940:8]
  wire  _T_301 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.TinyRocketConfig.fir 196963:6]
  wire  _T_309 = _T_20 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196972:8]
  wire  _T_310 = ~_T_309; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196973:8]
  wire  _T_320 = _T_17 & _T_32; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 196987:8]
  wire  _T_322 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.TinyRocketConfig.fir 196989:8]
  wire  _T_360 = _T_27 | _T_37; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197027:8]
  wire  _T_361 = _T_360 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197028:8]
  wire  _T_362 = _T_361 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197029:8]
  wire  _T_363 = _T_362 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197030:8]
  wire  _T_364 = _T_363 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197031:8]
  wire  _T_365 = _T_364 | _T_62; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197032:8]
  wire  _T_366 = _T_322 & _T_365; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 197033:8]
  wire  _T_368 = _T_320 | _T_366; // @[Parameters.scala 672:30 chipyard.TestHarness.TinyRocketConfig.fir 197035:8]
  wire  _T_370 = _T_368 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197037:8]
  wire  _T_371 = ~_T_370; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197038:8]
  wire  _T_378 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.TinyRocketConfig.fir 197057:8]
  wire  _T_380 = _T_378 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197059:8]
  wire  _T_381 = ~_T_380; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197060:8]
  wire  _T_382 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.TinyRocketConfig.fir 197065:8]
  wire  _T_384 = _T_382 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197067:8]
  wire  _T_385 = ~_T_384; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197068:8]
  wire  _T_390 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.TinyRocketConfig.fir 197082:6]
  wire  _T_441 = _T_27 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197134:8]
  wire  _T_442 = _T_441 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197135:8]
  wire  _T_443 = _T_442 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197136:8]
  wire  _T_444 = _T_443 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197137:8]
  wire  _T_445 = _T_444 | _T_62; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197138:8]
  wire  _T_446 = _T_322 & _T_445; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 197139:8]
  wire  _T_455 = _T_320 | _T_446; // @[Parameters.scala 672:30 chipyard.TestHarness.TinyRocketConfig.fir 197148:8]
  wire  _T_457 = _T_20 & _T_455; // @[Monitor.scala 115:71 chipyard.TestHarness.TinyRocketConfig.fir 197150:8]
  wire  _T_459 = _T_457 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197152:8]
  wire  _T_460 = ~_T_459; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197153:8]
  wire  _T_475 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.TinyRocketConfig.fir 197189:6]
  wire [3:0] _T_556 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.TinyRocketConfig.fir 197287:8]
  wire [3:0] _T_557 = io_in_a_bits_mask & _T_556; // @[Monitor.scala 127:31 chipyard.TestHarness.TinyRocketConfig.fir 197288:8]
  wire  _T_558 = _T_557 == 4'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.TinyRocketConfig.fir 197289:8]
  wire  _T_560 = _T_558 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197291:8]
  wire  _T_561 = ~_T_560; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197292:8]
  wire  _T_562 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.TinyRocketConfig.fir 197298:6]
  wire  _T_570 = io_in_a_bits_size <= 4'h2; // @[Parameters.scala 92:42 chipyard.TestHarness.TinyRocketConfig.fir 197307:8]
  wire  _T_609 = _T_63 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197346:8]
  wire  _T_610 = _T_609 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197347:8]
  wire  _T_611 = _T_610 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197348:8]
  wire  _T_612 = _T_611 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197349:8]
  wire  _T_613 = _T_612 | _T_62; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 197350:8]
  wire  _T_614 = _T_570 & _T_613; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 197351:8]
  wire  _T_624 = _T_20 & _T_614; // @[Monitor.scala 131:74 chipyard.TestHarness.TinyRocketConfig.fir 197361:8]
  wire  _T_626 = _T_624 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197363:8]
  wire  _T_627 = ~_T_626; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197364:8]
  wire  _T_634 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.TinyRocketConfig.fir 197383:8]
  wire  _T_636 = _T_634 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197385:8]
  wire  _T_637 = ~_T_636; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197386:8]
  wire  _T_642 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.TinyRocketConfig.fir 197400:6]
  wire  _T_714 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.TinyRocketConfig.fir 197485:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197487:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197488:8]
  wire  _T_722 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.TinyRocketConfig.fir 197502:6]
  wire  _T_784 = _T_20 & _T_320; // @[Monitor.scala 147:68 chipyard.TestHarness.TinyRocketConfig.fir 197565:8]
  wire  _T_786 = _T_784 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197567:8]
  wire  _T_787 = ~_T_786; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197568:8]
  wire  _T_794 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.TinyRocketConfig.fir 197587:8]
  wire  _T_796 = _T_794 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197589:8]
  wire  _T_797 = ~_T_796; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197590:8]
  wire  _T_806 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.TinyRocketConfig.fir 197614:6]
  wire  _T_808 = _T_806 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197616:6]
  wire  _T_809 = ~_T_808; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197617:6]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.TinyRocketConfig.fir 197622:6]
  wire  _T_810 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.TinyRocketConfig.fir 197627:6]
  wire  _T_812 = _source_ok_T_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197630:8]
  wire  _T_813 = ~_T_812; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197631:8]
  wire  _T_814 = io_in_d_bits_size >= 4'h2; // @[Monitor.scala 312:27 chipyard.TestHarness.TinyRocketConfig.fir 197636:8]
  wire  _T_816 = _T_814 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197638:8]
  wire  _T_817 = ~_T_816; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197639:8]
  wire  _T_818 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.TinyRocketConfig.fir 197644:8]
  wire  _T_820 = _T_818 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197646:8]
  wire  _T_821 = ~_T_820; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197647:8]
  wire  _T_822 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.TinyRocketConfig.fir 197652:8]
  wire  _T_824 = _T_822 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197654:8]
  wire  _T_825 = ~_T_824; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197655:8]
  wire  _T_826 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.TinyRocketConfig.fir 197660:8]
  wire  _T_828 = _T_826 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197662:8]
  wire  _T_829 = ~_T_828; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197663:8]
  wire  _T_830 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.TinyRocketConfig.fir 197669:6]
  wire  _T_841 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.TinyRocketConfig.fir 197693:8]
  wire  _T_843 = _T_841 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197695:8]
  wire  _T_844 = ~_T_843; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197696:8]
  wire  _T_845 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.TinyRocketConfig.fir 197701:8]
  wire  _T_847 = _T_845 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197703:8]
  wire  _T_848 = ~_T_847; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197704:8]
  wire  _T_858 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.TinyRocketConfig.fir 197727:6]
  wire  _T_878 = _T_826 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.TinyRocketConfig.fir 197768:8]
  wire  _T_880 = _T_878 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197770:8]
  wire  _T_881 = ~_T_880; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197771:8]
  wire  _T_887 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.TinyRocketConfig.fir 197786:6]
  wire  _T_904 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.TinyRocketConfig.fir 197821:6]
  wire  _T_922 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.TinyRocketConfig.fir 197857:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 197923:4]
  wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2]; // @[Edges.scala 219:59 chipyard.TestHarness.TinyRocketConfig.fir 197928:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.TinyRocketConfig.fir 197930:4]
  reg [9:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 197932:4]
  wire [9:0] a_first_counter1 = a_first_counter - 10'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 197934:4]
  wire  a_first = a_first_counter == 10'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 197935:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.TinyRocketConfig.fir 197946:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.TinyRocketConfig.fir 197947:4]
  reg [3:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.TinyRocketConfig.fir 197948:4]
  reg  source; // @[Monitor.scala 387:22 chipyard.TestHarness.TinyRocketConfig.fir 197949:4]
  reg [31:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.TinyRocketConfig.fir 197950:4]
  wire  _T_951 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.TinyRocketConfig.fir 197951:4]
  wire  _T_952 = io_in_a_valid & _T_951; // @[Monitor.scala 389:19 chipyard.TestHarness.TinyRocketConfig.fir 197952:4]
  wire  _T_953 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.TinyRocketConfig.fir 197954:6]
  wire  _T_955 = _T_953 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197956:6]
  wire  _T_956 = ~_T_955; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197957:6]
  wire  _T_957 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.TinyRocketConfig.fir 197962:6]
  wire  _T_959 = _T_957 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197964:6]
  wire  _T_960 = ~_T_959; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197965:6]
  wire  _T_961 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.TinyRocketConfig.fir 197970:6]
  wire  _T_963 = _T_961 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197972:6]
  wire  _T_964 = ~_T_963; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197973:6]
  wire  _T_965 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.TinyRocketConfig.fir 197978:6]
  wire  _T_967 = _T_965 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197980:6]
  wire  _T_968 = ~_T_967; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197981:6]
  wire  _T_969 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.TinyRocketConfig.fir 197986:6]
  wire  _T_971 = _T_969 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197988:6]
  wire  _T_972 = ~_T_971; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197989:6]
  wire  _T_974 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.TinyRocketConfig.fir 197996:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 198004:4]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 198006:4]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 198008:4]
  wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2]; // @[Edges.scala 219:59 chipyard.TestHarness.TinyRocketConfig.fir 198009:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.TinyRocketConfig.fir 198010:4]
  reg [9:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198012:4]
  wire [9:0] d_first_counter1 = d_first_counter - 10'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 198014:4]
  wire  d_first = d_first_counter == 10'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 198015:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.TinyRocketConfig.fir 198026:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.TinyRocketConfig.fir 198027:4]
  reg [3:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.TinyRocketConfig.fir 198028:4]
  reg  source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.TinyRocketConfig.fir 198029:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.TinyRocketConfig.fir 198030:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.TinyRocketConfig.fir 198031:4]
  wire  _T_975 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.TinyRocketConfig.fir 198032:4]
  wire  _T_976 = io_in_d_valid & _T_975; // @[Monitor.scala 541:19 chipyard.TestHarness.TinyRocketConfig.fir 198033:4]
  wire  _T_977 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.TinyRocketConfig.fir 198035:6]
  wire  _T_979 = _T_977 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198037:6]
  wire  _T_980 = ~_T_979; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198038:6]
  wire  _T_981 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.TinyRocketConfig.fir 198043:6]
  wire  _T_983 = _T_981 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198045:6]
  wire  _T_984 = ~_T_983; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198046:6]
  wire  _T_985 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.TinyRocketConfig.fir 198051:6]
  wire  _T_987 = _T_985 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198053:6]
  wire  _T_988 = ~_T_987; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198054:6]
  wire  _T_989 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.TinyRocketConfig.fir 198059:6]
  wire  _T_991 = _T_989 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198061:6]
  wire  _T_992 = ~_T_991; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198062:6]
  wire  _T_993 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.TinyRocketConfig.fir 198067:6]
  wire  _T_995 = _T_993 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198069:6]
  wire  _T_996 = ~_T_995; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198070:6]
  wire  _T_997 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.TinyRocketConfig.fir 198075:6]
  wire  _T_999 = _T_997 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198077:6]
  wire  _T_1000 = ~_T_999; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198078:6]
  wire  _T_1002 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.TinyRocketConfig.fir 198085:4]
  reg  inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 198094:4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 198095:4]
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 198096:4]
  reg [9:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198106:4]
  wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 198108:4]
  wire  a_first_1 = a_first_counter_1 == 10'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 198109:4]
  reg [9:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198128:4]
  wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 198130:4]
  wire  d_first_1 = d_first_counter_1 == 10'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 198131:4]
  wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.TinyRocketConfig.fir 198152:4]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.TinyRocketConfig.fir 198152:4]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.TinyRocketConfig.fir 198153:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.TinyRocketConfig.fir 198157:4]
  wire [15:0] _GEN_73 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.TinyRocketConfig.fir 198158:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.TinyRocketConfig.fir 198158:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.TinyRocketConfig.fir 198159:4]
  wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65 chipyard.TestHarness.TinyRocketConfig.fir 198163:4]
  wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.TinyRocketConfig.fir 198164:4]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.TinyRocketConfig.fir 198168:4]
  wire [15:0] _GEN_75 = {{8'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.TinyRocketConfig.fir 198169:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.TinyRocketConfig.fir 198169:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.TinyRocketConfig.fir 198170:4]
  wire  _T_1003 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.TinyRocketConfig.fir 198194:4]
  wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.TinyRocketConfig.fir 198197:6]
  wire [1:0] _GEN_15 = _T_1003 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.TinyRocketConfig.fir 198196:4 Monitor.scala 649:22 chipyard.TestHarness.TinyRocketConfig.fir 198198:6 chipyard.TestHarness.TinyRocketConfig.fir 198145:4]
  wire  _T_1006 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.TinyRocketConfig.fir 198201:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.TinyRocketConfig.fir 198206:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.TinyRocketConfig.fir 198207:6]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.TinyRocketConfig.fir 198209:6]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.TinyRocketConfig.fir 198210:6]
  wire [2:0] _GEN_77 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.TinyRocketConfig.fir 198212:6]
  wire [3:0] _a_opcodes_set_T = {{1'd0}, _GEN_77}; // @[Monitor.scala 656:79 chipyard.TestHarness.TinyRocketConfig.fir 198212:6]
  wire [3:0] a_opcodes_set_interm = _T_1006 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 198203:4 Monitor.scala 654:28 chipyard.TestHarness.TinyRocketConfig.fir 198208:6 chipyard.TestHarness.TinyRocketConfig.fir 198191:4]
  wire [18:0] _GEN_78 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.TinyRocketConfig.fir 198213:6]
  wire [18:0] _a_opcodes_set_T_1 = _GEN_78 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.TinyRocketConfig.fir 198213:6]
  wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 657:77 chipyard.TestHarness.TinyRocketConfig.fir 198215:6]
  wire [4:0] a_sizes_set_interm = _T_1006 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 198203:4 Monitor.scala 655:28 chipyard.TestHarness.TinyRocketConfig.fir 198211:6 chipyard.TestHarness.TinyRocketConfig.fir 198193:4]
  wire [19:0] _GEN_79 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.TinyRocketConfig.fir 198216:6]
  wire [19:0] _a_sizes_set_T_1 = _GEN_79 << _a_sizes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.TinyRocketConfig.fir 198216:6]
  wire  _T_1008 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.TinyRocketConfig.fir 198218:6]
  wire  _T_1010 = ~_T_1008; // @[Monitor.scala 658:17 chipyard.TestHarness.TinyRocketConfig.fir 198220:6]
  wire  _T_1012 = _T_1010 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 198222:6]
  wire  _T_1013 = ~_T_1012; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 198223:6]
  wire [1:0] _GEN_16 = _T_1006 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 198203:4 Monitor.scala 653:28 chipyard.TestHarness.TinyRocketConfig.fir 198205:6 chipyard.TestHarness.TinyRocketConfig.fir 198143:4]
  wire [18:0] _GEN_19 = _T_1006 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 198203:4 Monitor.scala 656:28 chipyard.TestHarness.TinyRocketConfig.fir 198214:6 chipyard.TestHarness.TinyRocketConfig.fir 198147:4]
  wire [19:0] _GEN_20 = _T_1006 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 198203:4 Monitor.scala 657:28 chipyard.TestHarness.TinyRocketConfig.fir 198217:6 chipyard.TestHarness.TinyRocketConfig.fir 198149:4]
  wire  _T_1014 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.TinyRocketConfig.fir 198238:4]
  wire  _T_1016 = ~_T_810; // @[Monitor.scala 671:74 chipyard.TestHarness.TinyRocketConfig.fir 198240:4]
  wire  _T_1017 = _T_1014 & _T_1016; // @[Monitor.scala 671:71 chipyard.TestHarness.TinyRocketConfig.fir 198241:4]
  wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.TinyRocketConfig.fir 198243:6]
  wire [1:0] _GEN_21 = _T_1017 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.TinyRocketConfig.fir 198242:4 Monitor.scala 672:22 chipyard.TestHarness.TinyRocketConfig.fir 198244:6 chipyard.TestHarness.TinyRocketConfig.fir 198232:4]
  wire  _T_1019 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.TinyRocketConfig.fir 198247:4]
  wire  _T_1022 = _T_1019 & _T_1016; // @[Monitor.scala 675:72 chipyard.TestHarness.TinyRocketConfig.fir 198250:4]
  wire [30:0] _GEN_81 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.TinyRocketConfig.fir 198259:6]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_81 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.TinyRocketConfig.fir 198259:6]
  wire [30:0] _GEN_82 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74 chipyard.TestHarness.TinyRocketConfig.fir 198266:6]
  wire [30:0] _d_sizes_clr_T_5 = _GEN_82 << _a_size_lookup_T; // @[Monitor.scala 678:74 chipyard.TestHarness.TinyRocketConfig.fir 198266:6]
  wire [1:0] _GEN_22 = _T_1022 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 198251:4 Monitor.scala 676:21 chipyard.TestHarness.TinyRocketConfig.fir 198253:6 chipyard.TestHarness.TinyRocketConfig.fir 198230:4]
  wire [30:0] _GEN_23 = _T_1022 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 198251:4 Monitor.scala 677:21 chipyard.TestHarness.TinyRocketConfig.fir 198260:6 chipyard.TestHarness.TinyRocketConfig.fir 198234:4]
  wire [30:0] _GEN_24 = _T_1022 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 198251:4 Monitor.scala 678:21 chipyard.TestHarness.TinyRocketConfig.fir 198267:6 chipyard.TestHarness.TinyRocketConfig.fir 198236:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.TinyRocketConfig.fir 198276:6]
  wire  same_cycle_resp = _T_1003 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.TinyRocketConfig.fir 198277:6]
  wire  _T_1027 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.TinyRocketConfig.fir 198278:6]
  wire  _T_1029 = _T_1027 | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.TinyRocketConfig.fir 198280:6]
  wire  _T_1031 = _T_1029 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198282:6]
  wire  _T_1032 = ~_T_1031; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198283:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8]
  wire  _T_1033 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 198289:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 198290:8 Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 198290:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 198290:8 Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 198290:8]
  wire  _T_1034 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 198290:8]
  wire  _T_1035 = _T_1033 | _T_1034; // @[Monitor.scala 685:77 chipyard.TestHarness.TinyRocketConfig.fir 198291:8]
  wire  _T_1037 = _T_1035 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198293:8]
  wire  _T_1038 = ~_T_1037; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198294:8]
  wire  _T_1039 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.TinyRocketConfig.fir 198299:8]
  wire  _T_1041 = _T_1039 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198301:8]
  wire  _T_1042 = ~_T_1041; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198302:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198150:4 Monitor.scala 634:21 chipyard.TestHarness.TinyRocketConfig.fir 198160:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8]
  wire  _T_1044 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 198310:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 198312:8 Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 198312:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 198312:8 Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 198312:8]
  wire  _T_1046 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 198312:8]
  wire  _T_1047 = _T_1044 | _T_1046; // @[Monitor.scala 689:72 chipyard.TestHarness.TinyRocketConfig.fir 198313:8]
  wire  _T_1049 = _T_1047 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198315:8]
  wire  _T_1050 = ~_T_1049; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198316:8]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198161:4 Monitor.scala 638:19 chipyard.TestHarness.TinyRocketConfig.fir 198171:4]
  wire [7:0] _GEN_83 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.TinyRocketConfig.fir 198321:8]
  wire  _T_1051 = _GEN_83 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.TinyRocketConfig.fir 198321:8]
  wire  _T_1053 = _T_1051 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198323:8]
  wire  _T_1054 = ~_T_1053; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198324:8]
  wire  _T_1056 = _T_1014 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.TinyRocketConfig.fir 198332:4]
  wire  _T_1057 = _T_1056 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.TinyRocketConfig.fir 198333:4]
  wire  _T_1059 = _T_1057 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.TinyRocketConfig.fir 198335:4]
  wire  _T_1061 = _T_1059 & _T_1016; // @[Monitor.scala 694:116 chipyard.TestHarness.TinyRocketConfig.fir 198337:4]
  wire  _T_1062 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.TinyRocketConfig.fir 198339:6]
  wire  _T_1063 = _T_1062 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.TinyRocketConfig.fir 198340:6]
  wire  _T_1065 = _T_1063 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198342:6]
  wire  _T_1066 = ~_T_1065; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198343:6]
  wire  a_set_wo_ready = _GEN_15[0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198144:4]
  wire  d_clr_wo_ready = _GEN_21[0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198231:4]
  wire  _T_1067 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.TinyRocketConfig.fir 198349:4]
  wire  _T_1068 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.TinyRocketConfig.fir 198350:4]
  wire  _T_1069 = ~_T_1068; // @[Monitor.scala 699:51 chipyard.TestHarness.TinyRocketConfig.fir 198351:4]
  wire  _T_1070 = _T_1067 | _T_1069; // @[Monitor.scala 699:48 chipyard.TestHarness.TinyRocketConfig.fir 198352:4]
  wire  _T_1072 = _T_1070 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198354:4]
  wire  _T_1073 = ~_T_1072; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198355:4]
  wire  a_set = _GEN_16[0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198142:4]
  wire  _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.TinyRocketConfig.fir 198360:4]
  wire  d_clr = _GEN_22[0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198229:4]
  wire  _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.TinyRocketConfig.fir 198361:4]
  wire  _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.TinyRocketConfig.fir 198362:4]
  wire [3:0] a_opcodes_set = _GEN_19[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198146:4]
  wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.TinyRocketConfig.fir 198364:4]
  wire [3:0] d_opcodes_clr = _GEN_23[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198233:4]
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.TinyRocketConfig.fir 198365:4]
  wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.TinyRocketConfig.fir 198366:4]
  wire [7:0] a_sizes_set = _GEN_20[7:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198148:4]
  wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.TinyRocketConfig.fir 198368:4]
  wire [7:0] d_sizes_clr = _GEN_24[7:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198235:4]
  wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56 chipyard.TestHarness.TinyRocketConfig.fir 198369:4]
  wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.TinyRocketConfig.fir 198370:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 198372:4]
  wire  _T_1074 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.TinyRocketConfig.fir 198375:4]
  wire  _T_1075 = ~_T_1074; // @[Monitor.scala 709:16 chipyard.TestHarness.TinyRocketConfig.fir 198376:4]
  wire  _T_1076 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.TinyRocketConfig.fir 198377:4]
  wire  _T_1077 = _T_1075 | _T_1076; // @[Monitor.scala 709:30 chipyard.TestHarness.TinyRocketConfig.fir 198378:4]
  wire  _T_1078 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.TinyRocketConfig.fir 198379:4]
  wire  _T_1079 = _T_1077 | _T_1078; // @[Monitor.scala 709:47 chipyard.TestHarness.TinyRocketConfig.fir 198380:4]
  wire  _T_1081 = _T_1079 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 198382:4]
  wire  _T_1082 = ~_T_1081; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 198383:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.TinyRocketConfig.fir 198389:4]
  wire  _T_1085 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.TinyRocketConfig.fir 198393:4]
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 198399:4]
  reg [9:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198434:4]
  wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 198436:4]
  wire  d_first_2 = d_first_counter_2 == 10'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 198437:4]
  wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.TinyRocketConfig.fir 198470:4]
  wire [15:0] _GEN_87 = {{8'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.TinyRocketConfig.fir 198475:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_87 & _a_size_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.TinyRocketConfig.fir 198475:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.TinyRocketConfig.fir 198476:4]
  wire  _T_1103 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.TinyRocketConfig.fir 198554:4]
  wire  _T_1105 = _T_1103 & _T_810; // @[Monitor.scala 779:71 chipyard.TestHarness.TinyRocketConfig.fir 198556:4]
  wire  _T_1107 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.TinyRocketConfig.fir 198562:4]
  wire  _T_1109 = _T_1107 & _T_810; // @[Monitor.scala 783:72 chipyard.TestHarness.TinyRocketConfig.fir 198564:4]
  wire [30:0] _GEN_69 = _T_1109 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.TinyRocketConfig.fir 198565:4 Monitor.scala 786:21 chipyard.TestHarness.TinyRocketConfig.fir 198581:6 chipyard.TestHarness.TinyRocketConfig.fir 198552:4]
  wire  _T_1113 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.TinyRocketConfig.fir 198600:6]
  wire  _T_1117 = _T_1113 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198604:6]
  wire  _T_1118 = ~_T_1117; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198605:6]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198458:4 Monitor.scala 747:21 chipyard.TestHarness.TinyRocketConfig.fir 198477:4]
  wire  _T_1123 = _GEN_83 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.TinyRocketConfig.fir 198623:8]
  wire  _T_1125 = _T_1123 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198625:8]
  wire  _T_1126 = ~_T_1125; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198626:8]
  wire [7:0] d_sizes_clr_1 = _GEN_69[7:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 198551:4]
  wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58 chipyard.TestHarness.TinyRocketConfig.fir 198676:4]
  wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.TinyRocketConfig.fir 198677:4]
  wire  _GEN_93 = io_in_a_valid & _T_15; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196668:10]
  wire  _GEN_109 = io_in_a_valid & _T_156; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196843:10]
  wire  _GEN_127 = io_in_a_valid & _T_301; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196975:10]
  wire  _GEN_141 = io_in_a_valid & _T_390; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197155:10]
  wire  _GEN_151 = io_in_a_valid & _T_475; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197262:10]
  wire  _GEN_161 = io_in_a_valid & _T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197366:10]
  wire  _GEN_171 = io_in_a_valid & _T_642; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197468:10]
  wire  _GEN_181 = io_in_a_valid & _T_722; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197570:10]
  wire  _GEN_193 = io_in_d_valid & _T_810; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197633:10]
  wire  _GEN_203 = io_in_d_valid & _T_830; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197675:10]
  wire  _GEN_215 = io_in_d_valid & _T_858; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197733:10]
  wire  _GEN_227 = io_in_d_valid & _T_887; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197792:10]
  wire  _GEN_233 = io_in_d_valid & _T_904; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197827:10]
  wire  _GEN_239 = io_in_d_valid & _T_922; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197863:10]
  wire  _GEN_245 = _T_1017 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198296:10]
  wire  _GEN_250 = _T_1017 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198318:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 198373:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 198680:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 197932:4]
      a_first_counter <= 10'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 197932:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 197942:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 197943:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 197931:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 10'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_974) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 197997:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.TinyRocketConfig.fir 197998:6]
    end
    if (_T_974) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 197997:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.TinyRocketConfig.fir 197999:6]
    end
    if (_T_974) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 197997:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.TinyRocketConfig.fir 198000:6]
    end
    if (_T_974) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 197997:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.TinyRocketConfig.fir 198001:6]
    end
    if (_T_974) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 197997:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.TinyRocketConfig.fir 198002:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198012:4]
      d_first_counter <= 10'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198012:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 198022:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 198023:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 198011:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 10'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 198086:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.TinyRocketConfig.fir 198087:6]
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 198086:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.TinyRocketConfig.fir 198088:6]
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 198086:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.TinyRocketConfig.fir 198089:6]
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 198086:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.TinyRocketConfig.fir 198090:6]
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 198086:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.TinyRocketConfig.fir 198091:6]
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 198086:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.TinyRocketConfig.fir 198092:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 198094:4]
      inflight <= 1'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 198094:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.TinyRocketConfig.fir 198363:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 198095:4]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 198095:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.TinyRocketConfig.fir 198367:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 198096:4]
      inflight_sizes <= 8'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 198096:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.TinyRocketConfig.fir 198371:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198106:4]
      a_first_counter_1 <= 10'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198106:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 198116:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 198117:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 197931:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 10'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198128:4]
      d_first_counter_1 <= 10'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198128:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 198138:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 198139:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 198011:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 10'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 198372:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 198372:4]
    end else if (_T_1085) begin // @[Monitor.scala 712:47 chipyard.TestHarness.TinyRocketConfig.fir 198394:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.TinyRocketConfig.fir 198395:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.TinyRocketConfig.fir 198390:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 198399:4]
      inflight_sizes_1 <= 8'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 198399:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.TinyRocketConfig.fir 198678:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198434:4]
      d_first_counter_2 <= 10'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 198434:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 198444:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 198445:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 198011:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 10'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_15 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196668:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_75) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196669:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196729:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_75) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196730:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_135) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196736:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_135) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196737:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_139) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196744:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_139) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196745:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196751:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196752:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_146) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196759:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_146) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196760:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_151) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196768:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_151) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196769:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_155) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196776:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_155) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196777:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_156 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196843:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_75) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196844:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196904:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_75) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196905:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_135) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196911:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_135) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196912:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_139) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196919:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_139) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196920:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196926:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196927:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_146) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196934:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_146) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196935:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_291) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196942:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_291) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196943:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_151) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196951:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_151) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196952:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_155) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196959:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_155) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196960:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_301 & _T_310) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196975:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_310) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 196976:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_371) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197040:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_371) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197041:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_135) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197047:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_135) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197048:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197054:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197055:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_381) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197062:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_381) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197063:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_385) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197070:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_385) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197071:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_155) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197078:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_155) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197079:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & _T_460) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197155:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_460) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197156:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_135) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197162:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_135) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197163:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197169:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197170:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_381) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197177:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_381) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197178:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_385) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197185:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_385) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197186:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_475 & _T_460) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197262:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_460) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197263:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_135) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197269:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_135) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197270:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197276:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197277:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_381) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197284:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_381) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197285:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_561) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197294:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_561) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197295:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_562 & _T_627) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197366:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_627) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197367:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_135) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197373:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_135) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197374:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197380:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197381:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_637) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197388:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_637) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197389:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_385) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197396:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_385) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197397:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_642 & _T_627) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197468:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_627) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197469:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_135) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197475:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_135) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197476:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197482:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197483:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197490:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_717) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197491:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_385) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197498:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_385) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197499:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_722 & _T_787) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197570:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_787) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197571:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_135) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197577:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_135) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197578:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197584:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197585:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_797) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197592:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_797) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197593:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_385) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197600:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_385) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197601:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_155) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197608:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_155) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197609:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_809) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197619:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_809) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197620:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_810 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197633:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197634:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_817) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197641:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_817) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197642:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_821) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197649:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_821) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197650:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_825) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197657:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_825) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197658:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_829) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197665:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_829) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197666:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_830 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197675:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197676:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197682:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_75) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197683:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_817) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197690:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_817) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197691:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_844) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197698:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_844) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197699:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_848) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197706:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_848) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197707:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_825) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197714:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_825) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197715:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_858 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197733:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197734:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197740:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_75) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197741:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_817) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197748:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_817) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197749:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_844) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197756:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_844) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197757:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_848) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197764:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_848) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197765:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_881) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197773:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_881) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197774:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_887 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197792:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197793:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_821) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197800:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_821) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197801:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_825) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197808:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_825) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197809:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_904 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197827:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197828:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_821) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197835:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_821) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197836:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_881) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197844:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_881) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197845:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_922 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197863:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_239 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197864:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_239 & _T_821) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197871:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_239 & _T_821) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197872:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_239 & _T_825) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197879:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_239 & _T_825) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 197880:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_952 & _T_956) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197959:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_952 & _T_956) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197960:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_952 & _T_960) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197967:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_952 & _T_960) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197968:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_952 & _T_964) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197975:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_952 & _T_964) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197976:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_952 & _T_968) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197983:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_952 & _T_968) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197984:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_952 & _T_972) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197991:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_952 & _T_972) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 197992:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_980) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198040:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_980) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198041:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_984) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198048:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_984) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198049:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_988) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198056:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_988) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198057:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_992) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198064:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_992) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198065:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_996) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198072:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_996) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198073:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_1000) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198080:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_1000) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198081:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1006 & _T_1013) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 198225:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1006 & _T_1013) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 198226:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1017 & _T_1032) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198285:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1017 & _T_1032) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198286:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1017 & same_cycle_resp & _T_1038) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198296:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_245 & _T_1038) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198297:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_245 & _T_1042) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198304:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_245 & _T_1042) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198305:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1017 & ~same_cycle_resp & _T_1050) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198318:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_250 & _T_1050) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198319:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_250 & _T_1054) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198326:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_250 & _T_1054) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198327:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1061 & _T_1066) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198345:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1061 & _T_1066) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198346:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1073) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 6 (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198357:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1073) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198358:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1082) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 198385:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1082) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 198386:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1105 & _T_1118) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198607:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1105 & _T_1118) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198608:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1105 & _T_1126) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198628:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1105 & _T_1126) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 198629:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inflight_opcodes = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  inflight_sizes = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[9:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[9:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_20[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLSerdesser_1_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 198891:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 198892:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 198893:4]
  output        auto_manager_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input         auto_manager_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [2:0]  auto_manager_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [2:0]  auto_manager_in_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [3:0]  auto_manager_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input         auto_manager_in_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [31:0] auto_manager_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [3:0]  auto_manager_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [31:0] auto_manager_in_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input         auto_manager_in_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input         auto_manager_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output        auto_manager_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [2:0]  auto_manager_in_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [1:0]  auto_manager_in_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [3:0]  auto_manager_in_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output        auto_manager_in_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output        auto_manager_in_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output        auto_manager_in_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [31:0] auto_manager_in_d_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output        auto_manager_in_d_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input         auto_client_out_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output        auto_client_out_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [2:0]  auto_client_out_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [2:0]  auto_client_out_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [2:0]  auto_client_out_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [1:0]  auto_client_out_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [28:0] auto_client_out_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [3:0]  auto_client_out_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output [31:0] auto_client_out_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output        auto_client_out_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output        auto_client_out_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input         auto_client_out_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [2:0]  auto_client_out_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [1:0]  auto_client_out_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [2:0]  auto_client_out_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [1:0]  auto_client_out_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input         auto_client_out_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input         auto_client_out_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input  [31:0] auto_client_out_d_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  input         auto_client_out_d_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 198894:4]
  output        io_ser_in_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 198895:4]
  input         io_ser_in_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 198895:4]
  input  [3:0]  io_ser_in_bits, // @[chipyard.TestHarness.TinyRocketConfig.fir 198895:4]
  input         io_ser_out_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 198895:4]
  output        io_ser_out_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 198895:4]
  output [3:0]  io_ser_out_bits // @[chipyard.TestHarness.TinyRocketConfig.fir 198895:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
  wire  outArb_clock; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_reset; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_in_1_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_in_1_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [2:0] outArb_io_in_1_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [2:0] outArb_io_in_1_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [3:0] outArb_io_in_1_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [1:0] outArb_io_in_1_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [31:0] outArb_io_in_1_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_in_1_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [3:0] outArb_io_in_1_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_in_1_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_in_4_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_in_4_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [2:0] outArb_io_in_4_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [2:0] outArb_io_in_4_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [3:0] outArb_io_in_4_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [1:0] outArb_io_in_4_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [31:0] outArb_io_in_4_bits_address; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [31:0] outArb_io_in_4_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_in_4_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [3:0] outArb_io_in_4_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_in_4_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_out_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_out_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [2:0] outArb_io_out_bits_chanId; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [2:0] outArb_io_out_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [2:0] outArb_io_out_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [3:0] outArb_io_out_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [1:0] outArb_io_out_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [31:0] outArb_io_out_bits_address; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [31:0] outArb_io_out_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_out_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire [3:0] outArb_io_out_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outArb_io_out_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
  wire  outSer_clock; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire  outSer_reset; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire  outSer_io_in_ready; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire  outSer_io_in_valid; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire [2:0] outSer_io_in_bits_chanId; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire [2:0] outSer_io_in_bits_opcode; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire [2:0] outSer_io_in_bits_param; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire [3:0] outSer_io_in_bits_size; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire [1:0] outSer_io_in_bits_source; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire [31:0] outSer_io_in_bits_address; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire [31:0] outSer_io_in_bits_data; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire  outSer_io_in_bits_corrupt; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire [3:0] outSer_io_in_bits_union; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire  outSer_io_in_bits_last; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire  outSer_io_out_ready; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire  outSer_io_out_valid; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire [3:0] outSer_io_out_bits; // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
  wire  inDes_clock; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire  inDes_reset; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire  inDes_io_in_ready; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire  inDes_io_in_valid; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire [3:0] inDes_io_in_bits; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire  inDes_io_out_ready; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire  inDes_io_out_valid; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire [2:0] inDes_io_out_bits_chanId; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire [2:0] inDes_io_out_bits_opcode; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire [2:0] inDes_io_out_bits_param; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire [3:0] inDes_io_out_bits_size; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire [1:0] inDes_io_out_bits_source; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire [31:0] inDes_io_out_bits_address; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire [31:0] inDes_io_out_bits_data; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire  inDes_io_out_bits_corrupt; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire [3:0] inDes_io_out_bits_union; // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
  wire [1:0] _merged_bits_merged_union_T_1 = {auto_client_out_d_bits_sink,auto_client_out_d_bits_denied}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 198994:4]
  wire  merged_1_ready = outArb_io_in_1_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.TinyRocketConfig.fir 198983:4 Serdes.scala 625:18 chipyard.TestHarness.TinyRocketConfig.fir 199179:4]
  wire  _merged_bits_last_T_1 = merged_1_ready & auto_client_out_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 199007:4]
  wire [12:0] _merged_bits_last_beats1_decode_T_1 = 13'h3f << auto_client_out_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 199009:4]
  wire [5:0] _merged_bits_last_beats1_decode_T_3 = ~_merged_bits_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 199011:4]
  wire [3:0] merged_bits_last_beats1_decode = _merged_bits_last_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59 chipyard.TestHarness.TinyRocketConfig.fir 199012:4]
  wire  merged_bits_last_beats1_opdata = auto_client_out_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.TinyRocketConfig.fir 199013:4]
  wire [3:0] merged_bits_last_beats1 = merged_bits_last_beats1_opdata ? merged_bits_last_beats1_decode : 4'h0; // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 199014:4]
  reg [3:0] merged_bits_last_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 199015:4]
  wire [3:0] merged_bits_last_counter1_1 = merged_bits_last_counter_1 - 4'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 199017:4]
  wire  merged_bits_last_first_1 = merged_bits_last_counter_1 == 4'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 199018:4]
  wire  _merged_bits_last_last_T_2 = merged_bits_last_counter_1 == 4'h1; // @[Edges.scala 231:25 chipyard.TestHarness.TinyRocketConfig.fir 199019:4]
  wire  _merged_bits_last_last_T_3 = merged_bits_last_beats1 == 4'h0; // @[Edges.scala 231:47 chipyard.TestHarness.TinyRocketConfig.fir 199020:4]
  wire  merged_4_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.TinyRocketConfig.fir 199126:4 Serdes.scala 625:18 chipyard.TestHarness.TinyRocketConfig.fir 199188:4]
  wire  _merged_bits_last_T_4 = merged_4_ready & auto_manager_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 199149:4]
  wire [20:0] _merged_bits_last_beats1_decode_T_13 = 21'h3f << auto_manager_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 199151:4]
  wire [5:0] _merged_bits_last_beats1_decode_T_15 = ~_merged_bits_last_beats1_decode_T_13[5:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 199153:4]
  wire [3:0] merged_bits_last_beats1_decode_3 = _merged_bits_last_beats1_decode_T_15[5:2]; // @[Edges.scala 219:59 chipyard.TestHarness.TinyRocketConfig.fir 199154:4]
  wire  merged_bits_last_beats1_opdata_3 = ~auto_manager_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.TinyRocketConfig.fir 199156:4]
  wire [3:0] merged_bits_last_beats1_3 = merged_bits_last_beats1_opdata_3 ? merged_bits_last_beats1_decode_3 : 4'h0; // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 199157:4]
  reg [3:0] merged_bits_last_counter_4; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 199158:4]
  wire [3:0] merged_bits_last_counter1_4 = merged_bits_last_counter_4 - 4'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 199160:4]
  wire  merged_bits_last_first_4 = merged_bits_last_counter_4 == 4'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 199161:4]
  wire  _merged_bits_last_last_T_8 = merged_bits_last_counter_4 == 4'h1; // @[Edges.scala 231:25 chipyard.TestHarness.TinyRocketConfig.fir 199162:4]
  wire  _merged_bits_last_last_T_9 = merged_bits_last_beats1_3 == 4'h0; // @[Edges.scala 231:47 chipyard.TestHarness.TinyRocketConfig.fir 199163:4]
  wire  _bundleOut_0_a_valid_T = inDes_io_out_bits_chanId == 3'h0; // @[Serdes.scala 236:37 chipyard.TestHarness.TinyRocketConfig.fir 199201:4]
  wire  _bundleIn_0_d_valid_T = inDes_io_out_bits_chanId == 3'h3; // @[Serdes.scala 239:37 chipyard.TestHarness.TinyRocketConfig.fir 199267:4]
  wire [3:0] _bundleIn_0_d_bits_d_sink_T = {{1'd0}, inDes_io_out_bits_union[3:1]}; // @[Serdes.scala 468:31 chipyard.TestHarness.TinyRocketConfig.fir 199277:4]
  wire  _inDes_io_out_ready_T = 3'h0 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.TinyRocketConfig.fir 199306:4]
  wire  _inDes_io_out_ready_T_1 = _inDes_io_out_ready_T & auto_client_out_a_ready; // @[Mux.scala 80:57 chipyard.TestHarness.TinyRocketConfig.fir 199307:4]
  wire  _inDes_io_out_ready_T_2 = 3'h1 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.TinyRocketConfig.fir 199308:4]
  wire  _inDes_io_out_ready_T_3 = _inDes_io_out_ready_T_2 ? 1'h0 : _inDes_io_out_ready_T_1; // @[Mux.scala 80:57 chipyard.TestHarness.TinyRocketConfig.fir 199309:4]
  wire  _inDes_io_out_ready_T_4 = 3'h2 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.TinyRocketConfig.fir 199310:4]
  wire  _inDes_io_out_ready_T_5 = _inDes_io_out_ready_T_4 ? 1'h0 : _inDes_io_out_ready_T_3; // @[Mux.scala 80:57 chipyard.TestHarness.TinyRocketConfig.fir 199311:4]
  wire  _inDes_io_out_ready_T_6 = 3'h3 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.TinyRocketConfig.fir 199312:4]
  wire  _inDes_io_out_ready_T_7 = _inDes_io_out_ready_T_6 ? auto_manager_in_d_ready : _inDes_io_out_ready_T_5; // @[Mux.scala 80:57 chipyard.TestHarness.TinyRocketConfig.fir 199313:4]
  wire  _inDes_io_out_ready_T_8 = 3'h4 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.TinyRocketConfig.fir 199314:4]
  TLMonitor_41_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 198905:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  HellaPeekingArbiter_inTestHarness outArb ( // @[Serdes.scala 622:24 chipyard.TestHarness.TinyRocketConfig.fir 198936:4]
    .clock(outArb_clock),
    .reset(outArb_reset),
    .io_in_1_ready(outArb_io_in_1_ready),
    .io_in_1_valid(outArb_io_in_1_valid),
    .io_in_1_bits_opcode(outArb_io_in_1_bits_opcode),
    .io_in_1_bits_param(outArb_io_in_1_bits_param),
    .io_in_1_bits_size(outArb_io_in_1_bits_size),
    .io_in_1_bits_source(outArb_io_in_1_bits_source),
    .io_in_1_bits_data(outArb_io_in_1_bits_data),
    .io_in_1_bits_corrupt(outArb_io_in_1_bits_corrupt),
    .io_in_1_bits_union(outArb_io_in_1_bits_union),
    .io_in_1_bits_last(outArb_io_in_1_bits_last),
    .io_in_4_ready(outArb_io_in_4_ready),
    .io_in_4_valid(outArb_io_in_4_valid),
    .io_in_4_bits_opcode(outArb_io_in_4_bits_opcode),
    .io_in_4_bits_param(outArb_io_in_4_bits_param),
    .io_in_4_bits_size(outArb_io_in_4_bits_size),
    .io_in_4_bits_source(outArb_io_in_4_bits_source),
    .io_in_4_bits_address(outArb_io_in_4_bits_address),
    .io_in_4_bits_data(outArb_io_in_4_bits_data),
    .io_in_4_bits_corrupt(outArb_io_in_4_bits_corrupt),
    .io_in_4_bits_union(outArb_io_in_4_bits_union),
    .io_in_4_bits_last(outArb_io_in_4_bits_last),
    .io_out_ready(outArb_io_out_ready),
    .io_out_valid(outArb_io_out_valid),
    .io_out_bits_chanId(outArb_io_out_bits_chanId),
    .io_out_bits_opcode(outArb_io_out_bits_opcode),
    .io_out_bits_param(outArb_io_out_bits_param),
    .io_out_bits_size(outArb_io_out_bits_size),
    .io_out_bits_source(outArb_io_out_bits_source),
    .io_out_bits_address(outArb_io_out_bits_address),
    .io_out_bits_data(outArb_io_out_bits_data),
    .io_out_bits_corrupt(outArb_io_out_bits_corrupt),
    .io_out_bits_union(outArb_io_out_bits_union),
    .io_out_bits_last(outArb_io_out_bits_last)
  );
  GenericSerializer_inTestHarness outSer ( // @[Serdes.scala 624:24 chipyard.TestHarness.TinyRocketConfig.fir 198939:4]
    .clock(outSer_clock),
    .reset(outSer_reset),
    .io_in_ready(outSer_io_in_ready),
    .io_in_valid(outSer_io_in_valid),
    .io_in_bits_chanId(outSer_io_in_bits_chanId),
    .io_in_bits_opcode(outSer_io_in_bits_opcode),
    .io_in_bits_param(outSer_io_in_bits_param),
    .io_in_bits_size(outSer_io_in_bits_size),
    .io_in_bits_source(outSer_io_in_bits_source),
    .io_in_bits_address(outSer_io_in_bits_address),
    .io_in_bits_data(outSer_io_in_bits_data),
    .io_in_bits_corrupt(outSer_io_in_bits_corrupt),
    .io_in_bits_union(outSer_io_in_bits_union),
    .io_in_bits_last(outSer_io_in_bits_last),
    .io_out_ready(outSer_io_out_ready),
    .io_out_valid(outSer_io_out_valid),
    .io_out_bits(outSer_io_out_bits)
  );
  GenericDeserializer_inTestHarness inDes ( // @[Serdes.scala 629:23 chipyard.TestHarness.TinyRocketConfig.fir 199195:4]
    .clock(inDes_clock),
    .reset(inDes_reset),
    .io_in_ready(inDes_io_in_ready),
    .io_in_valid(inDes_io_in_valid),
    .io_in_bits(inDes_io_in_bits),
    .io_out_ready(inDes_io_out_ready),
    .io_out_valid(inDes_io_out_valid),
    .io_out_bits_chanId(inDes_io_out_bits_chanId),
    .io_out_bits_opcode(inDes_io_out_bits_opcode),
    .io_out_bits_param(inDes_io_out_bits_param),
    .io_out_bits_size(inDes_io_out_bits_size),
    .io_out_bits_source(inDes_io_out_bits_source),
    .io_out_bits_address(inDes_io_out_bits_address),
    .io_out_bits_data(inDes_io_out_bits_data),
    .io_out_bits_corrupt(inDes_io_out_bits_corrupt),
    .io_out_bits_union(inDes_io_out_bits_union)
  );
  assign auto_manager_in_a_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.TinyRocketConfig.fir 199126:4 Serdes.scala 625:18 chipyard.TestHarness.TinyRocketConfig.fir 199188:4]
  assign auto_manager_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 637:46 chipyard.TestHarness.TinyRocketConfig.fir 199268:4]
  assign auto_manager_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 461:15 chipyard.TestHarness.TinyRocketConfig.fir 199271:4]
  assign auto_manager_in_d_bits_param = inDes_io_out_bits_param[1:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 462:15 chipyard.TestHarness.TinyRocketConfig.fir 199272:4]
  assign auto_manager_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 463:15 chipyard.TestHarness.TinyRocketConfig.fir 199273:4]
  assign auto_manager_in_d_bits_source = inDes_io_out_bits_source[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 464:15 chipyard.TestHarness.TinyRocketConfig.fir 199274:4]
  assign auto_manager_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 468:17 chipyard.TestHarness.TinyRocketConfig.fir 199278:4]
  assign auto_manager_in_d_bits_denied = inDes_io_out_bits_union[0]; // @[Serdes.scala 469:30 chipyard.TestHarness.TinyRocketConfig.fir 199279:4]
  assign auto_manager_in_d_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 465:15 chipyard.TestHarness.TinyRocketConfig.fir 199275:4]
  assign auto_manager_in_d_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 467:17 chipyard.TestHarness.TinyRocketConfig.fir 199276:4]
  assign auto_client_out_a_valid = inDes_io_out_valid & _bundleOut_0_a_valid_T; // @[Serdes.scala 631:45 chipyard.TestHarness.TinyRocketConfig.fir 199202:4]
  assign auto_client_out_a_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 374:17 chipyard.TestHarness.TinyRocketConfig.fir 199204:4 Serdes.scala 375:15 chipyard.TestHarness.TinyRocketConfig.fir 199205:4]
  assign auto_client_out_a_bits_param = inDes_io_out_bits_param; // @[Serdes.scala 374:17 chipyard.TestHarness.TinyRocketConfig.fir 199204:4 Serdes.scala 376:15 chipyard.TestHarness.TinyRocketConfig.fir 199206:4]
  assign auto_client_out_a_bits_size = inDes_io_out_bits_size[2:0]; // @[Serdes.scala 374:17 chipyard.TestHarness.TinyRocketConfig.fir 199204:4 Serdes.scala 377:15 chipyard.TestHarness.TinyRocketConfig.fir 199207:4]
  assign auto_client_out_a_bits_source = inDes_io_out_bits_source; // @[Serdes.scala 374:17 chipyard.TestHarness.TinyRocketConfig.fir 199204:4 Serdes.scala 378:15 chipyard.TestHarness.TinyRocketConfig.fir 199208:4]
  assign auto_client_out_a_bits_address = inDes_io_out_bits_address[28:0]; // @[Serdes.scala 374:17 chipyard.TestHarness.TinyRocketConfig.fir 199204:4 Serdes.scala 379:15 chipyard.TestHarness.TinyRocketConfig.fir 199209:4]
  assign auto_client_out_a_bits_mask = inDes_io_out_bits_union; // @[Serdes.scala 374:17 chipyard.TestHarness.TinyRocketConfig.fir 199204:4 Serdes.scala 385:15 chipyard.TestHarness.TinyRocketConfig.fir 199212:4]
  assign auto_client_out_a_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 374:17 chipyard.TestHarness.TinyRocketConfig.fir 199204:4 Serdes.scala 380:15 chipyard.TestHarness.TinyRocketConfig.fir 199210:4]
  assign auto_client_out_a_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 374:17 chipyard.TestHarness.TinyRocketConfig.fir 199204:4 Serdes.scala 382:17 chipyard.TestHarness.TinyRocketConfig.fir 199211:4]
  assign auto_client_out_d_ready = outArb_io_in_1_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.TinyRocketConfig.fir 198983:4 Serdes.scala 625:18 chipyard.TestHarness.TinyRocketConfig.fir 199179:4]
  assign io_ser_in_ready = inDes_io_in_ready; // @[Serdes.scala 630:17 chipyard.TestHarness.TinyRocketConfig.fir 199200:4]
  assign io_ser_out_valid = outSer_io_out_valid; // @[Serdes.scala 627:16 chipyard.TestHarness.TinyRocketConfig.fir 199193:4]
  assign io_ser_out_bits = outSer_io_out_bits; // @[Serdes.scala 627:16 chipyard.TestHarness.TinyRocketConfig.fir 199192:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 198906:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 198907:4]
  assign monitor_io_in_a_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.TinyRocketConfig.fir 199126:4 Serdes.scala 625:18 chipyard.TestHarness.TinyRocketConfig.fir 199188:4]
  assign monitor_io_in_a_valid = auto_manager_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign monitor_io_in_a_bits_opcode = auto_manager_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign monitor_io_in_a_bits_param = auto_manager_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign monitor_io_in_a_bits_size = auto_manager_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign monitor_io_in_a_bits_source = auto_manager_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign monitor_io_in_a_bits_address = auto_manager_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign monitor_io_in_a_bits_mask = auto_manager_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign monitor_io_in_a_bits_corrupt = auto_manager_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign monitor_io_in_d_ready = auto_manager_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign monitor_io_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 637:46 chipyard.TestHarness.TinyRocketConfig.fir 199268:4]
  assign monitor_io_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 461:15 chipyard.TestHarness.TinyRocketConfig.fir 199271:4]
  assign monitor_io_in_d_bits_param = inDes_io_out_bits_param[1:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 462:15 chipyard.TestHarness.TinyRocketConfig.fir 199272:4]
  assign monitor_io_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 463:15 chipyard.TestHarness.TinyRocketConfig.fir 199273:4]
  assign monitor_io_in_d_bits_source = inDes_io_out_bits_source[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 464:15 chipyard.TestHarness.TinyRocketConfig.fir 199274:4]
  assign monitor_io_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 468:17 chipyard.TestHarness.TinyRocketConfig.fir 199278:4]
  assign monitor_io_in_d_bits_denied = inDes_io_out_bits_union[0]; // @[Serdes.scala 469:30 chipyard.TestHarness.TinyRocketConfig.fir 199279:4]
  assign monitor_io_in_d_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 460:17 chipyard.TestHarness.TinyRocketConfig.fir 199270:4 Serdes.scala 467:17 chipyard.TestHarness.TinyRocketConfig.fir 199276:4]
  assign outArb_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 198937:4]
  assign outArb_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 198938:4]
  assign outArb_io_in_1_valid = auto_client_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 198901:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 198928:4]
  assign outArb_io_in_1_bits_opcode = auto_client_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 198901:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 198928:4]
  assign outArb_io_in_1_bits_param = {{1'd0}, auto_client_out_d_bits_param}; // @[Serdes.scala 312:22 chipyard.TestHarness.TinyRocketConfig.fir 198985:4 Serdes.scala 315:20 chipyard.TestHarness.TinyRocketConfig.fir 198988:4]
  assign outArb_io_in_1_bits_size = {{1'd0}, auto_client_out_d_bits_size}; // @[Serdes.scala 312:22 chipyard.TestHarness.TinyRocketConfig.fir 198985:4 Serdes.scala 316:20 chipyard.TestHarness.TinyRocketConfig.fir 198989:4]
  assign outArb_io_in_1_bits_source = auto_client_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 198901:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 198928:4]
  assign outArb_io_in_1_bits_data = auto_client_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 198901:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 198928:4]
  assign outArb_io_in_1_bits_corrupt = auto_client_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 198901:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 198928:4]
  assign outArb_io_in_1_bits_union = {{2'd0}, _merged_bits_merged_union_T_1}; // @[Serdes.scala 312:22 chipyard.TestHarness.TinyRocketConfig.fir 198985:4 Serdes.scala 322:22 chipyard.TestHarness.TinyRocketConfig.fir 198995:4]
  assign outArb_io_in_1_bits_last = _merged_bits_last_last_T_2 | _merged_bits_last_last_T_3; // @[Edges.scala 231:37 chipyard.TestHarness.TinyRocketConfig.fir 199021:4]
  assign outArb_io_in_4_valid = auto_manager_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign outArb_io_in_4_bits_opcode = auto_manager_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign outArb_io_in_4_bits_param = auto_manager_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign outArb_io_in_4_bits_size = auto_manager_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign outArb_io_in_4_bits_source = {{1'd0}, auto_manager_in_a_bits_source}; // @[Serdes.scala 255:22 chipyard.TestHarness.TinyRocketConfig.fir 199128:4 Serdes.scala 260:20 chipyard.TestHarness.TinyRocketConfig.fir 199133:4]
  assign outArb_io_in_4_bits_address = auto_manager_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign outArb_io_in_4_bits_data = auto_manager_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign outArb_io_in_4_bits_corrupt = auto_manager_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign outArb_io_in_4_bits_union = auto_manager_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 198903:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 198929:4]
  assign outArb_io_in_4_bits_last = _merged_bits_last_last_T_8 | _merged_bits_last_last_T_9; // @[Edges.scala 231:37 chipyard.TestHarness.TinyRocketConfig.fir 199164:4]
  assign outArb_io_out_ready = outSer_io_in_ready; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199191:4]
  assign outSer_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 198940:4]
  assign outSer_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 198941:4]
  assign outSer_io_in_valid = outArb_io_out_valid; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199190:4]
  assign outSer_io_in_bits_chanId = outArb_io_out_bits_chanId; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199189:4]
  assign outSer_io_in_bits_opcode = outArb_io_out_bits_opcode; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199189:4]
  assign outSer_io_in_bits_param = outArb_io_out_bits_param; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199189:4]
  assign outSer_io_in_bits_size = outArb_io_out_bits_size; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199189:4]
  assign outSer_io_in_bits_source = outArb_io_out_bits_source; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199189:4]
  assign outSer_io_in_bits_address = outArb_io_out_bits_address; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199189:4]
  assign outSer_io_in_bits_data = outArb_io_out_bits_data; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199189:4]
  assign outSer_io_in_bits_corrupt = outArb_io_out_bits_corrupt; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199189:4]
  assign outSer_io_in_bits_union = outArb_io_out_bits_union; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199189:4]
  assign outSer_io_in_bits_last = outArb_io_out_bits_last; // @[Serdes.scala 626:18 chipyard.TestHarness.TinyRocketConfig.fir 199189:4]
  assign outSer_io_out_ready = io_ser_out_ready; // @[Serdes.scala 627:16 chipyard.TestHarness.TinyRocketConfig.fir 199194:4]
  assign inDes_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 199196:4]
  assign inDes_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 199197:4]
  assign inDes_io_in_valid = io_ser_in_valid; // @[Serdes.scala 630:17 chipyard.TestHarness.TinyRocketConfig.fir 199199:4]
  assign inDes_io_in_bits = io_ser_in_bits; // @[Serdes.scala 630:17 chipyard.TestHarness.TinyRocketConfig.fir 199198:4]
  assign inDes_io_out_ready = _inDes_io_out_ready_T_8 ? 1'h0 : _inDes_io_out_ready_T_7; // @[Mux.scala 80:57 chipyard.TestHarness.TinyRocketConfig.fir 199315:4]
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 199015:4]
      merged_bits_last_counter_1 <= 4'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 199015:4]
    end else if (_merged_bits_last_T_1) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 199025:4]
      if (merged_bits_last_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 199026:6]
        if (merged_bits_last_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 199014:4]
          merged_bits_last_counter_1 <= merged_bits_last_beats1_decode;
        end else begin
          merged_bits_last_counter_1 <= 4'h0;
        end
      end else begin
        merged_bits_last_counter_1 <= merged_bits_last_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 199158:4]
      merged_bits_last_counter_4 <= 4'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 199158:4]
    end else if (_merged_bits_last_T_4) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 199168:4]
      if (merged_bits_last_first_4) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 199169:6]
        if (merged_bits_last_beats1_opdata_3) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 199157:4]
          merged_bits_last_counter_4 <= merged_bits_last_beats1_decode_3;
        end else begin
          merged_bits_last_counter_4 <= 4'h0;
        end
      end else begin
        merged_bits_last_counter_4 <= merged_bits_last_counter1_4;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  merged_bits_last_counter_1 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  merged_bits_last_counter_4 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_42_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 199334:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 199335:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 199336:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input  [1:0]  io_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input  [6:0]  io_in_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input  [3:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input  [1:0]  io_in_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
  input  [6:0]  io_in_d_bits_source // @[chipyard.TestHarness.TinyRocketConfig.fir 199337:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [95:0] _RAND_10;
  reg [383:0] _RAND_11;
  reg [383:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [95:0] _RAND_16;
  reg [383:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 200797:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 201104:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 7'h5f; // @[Parameters.scala 57:20 chipyard.TestHarness.TinyRocketConfig.fir 199354:6]
  wire [4:0] _is_aligned_mask_T_1 = 5'h3 << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 199360:6]
  wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 199362:6]
  wire [28:0] _GEN_71 = {{27'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.TinyRocketConfig.fir 199363:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.TinyRocketConfig.fir 199363:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.TinyRocketConfig.fir 199364:6]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49 chipyard.TestHarness.TinyRocketConfig.fir 199366:6]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.TinyRocketConfig.fir 199367:6]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81 chipyard.TestHarness.TinyRocketConfig.fir 199369:6]
  wire  _mask_T = io_in_a_bits_size >= 2'h2; // @[Misc.scala 205:21 chipyard.TestHarness.TinyRocketConfig.fir 199370:6]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 199371:6]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 199372:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 199373:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 199375:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 199376:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 199378:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 199379:6]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 199380:6]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 199381:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 199382:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 199383:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 199384:6]
  wire  mask_lo_lo = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 199385:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 199386:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 199387:6]
  wire  mask_lo_hi = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 199388:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 199389:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 199390:6]
  wire  mask_hi_lo = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 199391:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 199392:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 199393:6]
  wire  mask_hi_hi = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 199394:6]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 199397:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.TinyRocketConfig.fir 199420:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 199436:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 199437:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 199439:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 199440:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199446:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199471:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199472:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199479:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199480:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199486:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199487:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.TinyRocketConfig.fir 199492:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199494:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199495:8]
  wire [3:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.TinyRocketConfig.fir 199500:8]
  wire  _T_74 = _T_73 == 4'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.TinyRocketConfig.fir 199501:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199503:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199504:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.TinyRocketConfig.fir 199509:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199511:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199512:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.TinyRocketConfig.fir 199518:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.TinyRocketConfig.fir 199598:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199600:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199601:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.TinyRocketConfig.fir 199624:6]
  wire  _T_164 = io_in_a_bits_size <= 2'h2; // @[Parameters.scala 92:42 chipyard.TestHarness.TinyRocketConfig.fir 199647:8]
  wire  _T_172 = _T_164 & _T_37; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 199655:8]
  wire  _T_175 = _T_172 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199658:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199659:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.TinyRocketConfig.fir 199678:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199680:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199681:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.TinyRocketConfig.fir 199686:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199688:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199689:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.TinyRocketConfig.fir 199703:6]
  wire  _T_218 = _source_ok_T_4 & _T_172; // @[Monitor.scala 115:71 chipyard.TestHarness.TinyRocketConfig.fir 199729:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199731:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199732:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.TinyRocketConfig.fir 199768:6]
  wire [3:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.TinyRocketConfig.fir 199824:8]
  wire [3:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.TinyRocketConfig.fir 199825:8]
  wire  _T_275 = _T_274 == 4'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.TinyRocketConfig.fir 199826:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199828:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199829:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.TinyRocketConfig.fir 199835:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.TinyRocketConfig.fir 199880:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199882:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199883:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.TinyRocketConfig.fir 199897:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.TinyRocketConfig.fir 199942:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199944:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199945:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.TinyRocketConfig.fir 199959:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.TinyRocketConfig.fir 200004:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200006:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200007:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.TinyRocketConfig.fir 200031:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200033:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200034:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 7'h5f; // @[Parameters.scala 57:20 chipyard.TestHarness.TinyRocketConfig.fir 200045:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.TinyRocketConfig.fir 200051:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200054:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200055:8]
  wire  _T_405 = io_in_d_bits_size >= 2'h2; // @[Monitor.scala 312:27 chipyard.TestHarness.TinyRocketConfig.fir 200060:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200062:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200063:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.TinyRocketConfig.fir 200093:6]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.TinyRocketConfig.fir 200151:6]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.TinyRocketConfig.fir 200210:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.TinyRocketConfig.fir 200245:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.TinyRocketConfig.fir 200281:6]
  wire  a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 200347:4]
  reg  a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200356:4]
  wire  a_first_counter1 = a_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 200358:4]
  wire  a_first = ~a_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 200359:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.TinyRocketConfig.fir 200370:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.TinyRocketConfig.fir 200371:4]
  reg [1:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.TinyRocketConfig.fir 200372:4]
  reg [6:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.TinyRocketConfig.fir 200373:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.TinyRocketConfig.fir 200374:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.TinyRocketConfig.fir 200375:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.TinyRocketConfig.fir 200376:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.TinyRocketConfig.fir 200378:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200380:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200381:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.TinyRocketConfig.fir 200386:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200388:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200389:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.TinyRocketConfig.fir 200394:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200396:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200397:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.TinyRocketConfig.fir 200402:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200404:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200405:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.TinyRocketConfig.fir 200410:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200412:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200413:6]
  wire  _T_565 = a_first_done & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.TinyRocketConfig.fir 200420:4]
  wire  d_first_done = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 200428:4]
  reg  d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200436:4]
  wire  d_first_counter1 = d_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 200438:4]
  wire  d_first = ~d_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 200439:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.TinyRocketConfig.fir 200450:4]
  reg [1:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.TinyRocketConfig.fir 200452:4]
  reg [6:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.TinyRocketConfig.fir 200453:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.TinyRocketConfig.fir 200456:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.TinyRocketConfig.fir 200457:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.TinyRocketConfig.fir 200459:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200461:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200462:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.TinyRocketConfig.fir 200475:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200477:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200478:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.TinyRocketConfig.fir 200483:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200485:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200486:6]
  wire  _T_593 = d_first_done & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.TinyRocketConfig.fir 200509:4]
  reg [95:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 200518:4]
  reg [383:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 200519:4]
  reg [383:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 200520:4]
  reg  a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200530:4]
  wire  a_first_counter1_1 = a_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 200532:4]
  wire  a_first_1 = ~a_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 200533:4]
  reg  d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200552:4]
  wire  d_first_counter1_1 = d_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 200554:4]
  wire  d_first_1 = ~d_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 200555:4]
  wire [8:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.TinyRocketConfig.fir 200576:4]
  wire [9:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.TinyRocketConfig.fir 200576:4]
  wire [383:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.TinyRocketConfig.fir 200577:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.TinyRocketConfig.fir 200581:4]
  wire [383:0] _GEN_73 = {{368'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.TinyRocketConfig.fir 200582:4]
  wire [383:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.TinyRocketConfig.fir 200582:4]
  wire [383:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[383:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.TinyRocketConfig.fir 200583:4]
  wire [383:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.TinyRocketConfig.fir 200588:4]
  wire [383:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.TinyRocketConfig.fir 200593:4]
  wire [383:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[383:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.TinyRocketConfig.fir 200594:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.TinyRocketConfig.fir 200618:4]
  wire [127:0] _a_set_wo_ready_T = 128'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.TinyRocketConfig.fir 200621:6]
  wire [127:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.TinyRocketConfig.fir 200620:4 Monitor.scala 649:22 chipyard.TestHarness.TinyRocketConfig.fir 200622:6 chipyard.TestHarness.TinyRocketConfig.fir 200569:4]
  wire  _T_597 = a_first_done & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.TinyRocketConfig.fir 200625:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.TinyRocketConfig.fir 200630:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.TinyRocketConfig.fir 200631:6]
  wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.TinyRocketConfig.fir 200633:6]
  wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.TinyRocketConfig.fir 200634:6]
  wire [8:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.TinyRocketConfig.fir 200636:6]
  wire [9:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.TinyRocketConfig.fir 200636:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 200627:4 Monitor.scala 654:28 chipyard.TestHarness.TinyRocketConfig.fir 200632:6 chipyard.TestHarness.TinyRocketConfig.fir 200615:4]
  wire [1026:0] _GEN_79 = {{1023'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.TinyRocketConfig.fir 200637:6]
  wire [1026:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.TinyRocketConfig.fir 200637:6]
  wire [2:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 3'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 200627:4 Monitor.scala 655:28 chipyard.TestHarness.TinyRocketConfig.fir 200635:6 chipyard.TestHarness.TinyRocketConfig.fir 200617:4]
  wire [1025:0] _GEN_81 = {{1023'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.TinyRocketConfig.fir 200640:6]
  wire [1025:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.TinyRocketConfig.fir 200640:6]
  wire [95:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.TinyRocketConfig.fir 200642:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.TinyRocketConfig.fir 200644:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200646:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200647:6]
  wire [127:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 200627:4 Monitor.scala 653:28 chipyard.TestHarness.TinyRocketConfig.fir 200629:6 chipyard.TestHarness.TinyRocketConfig.fir 200567:4]
  wire [1026:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 200627:4 Monitor.scala 656:28 chipyard.TestHarness.TinyRocketConfig.fir 200638:6 chipyard.TestHarness.TinyRocketConfig.fir 200571:4]
  wire [1025:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 1026'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 200627:4 Monitor.scala 657:28 chipyard.TestHarness.TinyRocketConfig.fir 200641:6 chipyard.TestHarness.TinyRocketConfig.fir 200573:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.TinyRocketConfig.fir 200662:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.TinyRocketConfig.fir 200664:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.TinyRocketConfig.fir 200665:4]
  wire [127:0] _d_clr_wo_ready_T = 128'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.TinyRocketConfig.fir 200667:6]
  wire [127:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.TinyRocketConfig.fir 200666:4 Monitor.scala 672:22 chipyard.TestHarness.TinyRocketConfig.fir 200668:6 chipyard.TestHarness.TinyRocketConfig.fir 200656:4]
  wire  _T_610 = d_first_done & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.TinyRocketConfig.fir 200671:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.TinyRocketConfig.fir 200674:4]
  wire [1038:0] _GEN_83 = {{1023'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.TinyRocketConfig.fir 200683:6]
  wire [1038:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.TinyRocketConfig.fir 200683:6]
  wire [127:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 200675:4 Monitor.scala 676:21 chipyard.TestHarness.TinyRocketConfig.fir 200677:6 chipyard.TestHarness.TinyRocketConfig.fir 200654:4]
  wire [1038:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 200675:4 Monitor.scala 677:21 chipyard.TestHarness.TinyRocketConfig.fir 200684:6 chipyard.TestHarness.TinyRocketConfig.fir 200658:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.TinyRocketConfig.fir 200700:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.TinyRocketConfig.fir 200701:6]
  wire [95:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.TinyRocketConfig.fir 200702:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.TinyRocketConfig.fir 200704:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200706:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200707:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 200713:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 200714:8 Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 200714:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 200714:8 Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 200714:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 200714:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.TinyRocketConfig.fir 200715:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200717:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200718:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.TinyRocketConfig.fir 200723:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200725:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200726:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200574:4 Monitor.scala 634:21 chipyard.TestHarness.TinyRocketConfig.fir 200584:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 200734:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 200736:8 Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 200736:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 200736:8 Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 200736:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 200736:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.TinyRocketConfig.fir 200737:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200739:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200740:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200585:4 Monitor.scala 638:19 chipyard.TestHarness.TinyRocketConfig.fir 200595:4]
  wire [3:0] _GEN_86 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.TinyRocketConfig.fir 200745:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.TinyRocketConfig.fir 200745:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200747:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200748:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.TinyRocketConfig.fir 200756:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.TinyRocketConfig.fir 200757:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.TinyRocketConfig.fir 200759:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.TinyRocketConfig.fir 200761:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.TinyRocketConfig.fir 200763:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.TinyRocketConfig.fir 200764:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200766:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200767:6]
  wire [95:0] a_set_wo_ready = _GEN_15[95:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200568:4]
  wire [95:0] d_clr_wo_ready = _GEN_21[95:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200655:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.TinyRocketConfig.fir 200773:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.TinyRocketConfig.fir 200774:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.TinyRocketConfig.fir 200775:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.TinyRocketConfig.fir 200776:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200778:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200779:4]
  wire [95:0] a_set = _GEN_16[95:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200566:4]
  wire [95:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.TinyRocketConfig.fir 200784:4]
  wire [95:0] d_clr = _GEN_22[95:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200653:4]
  wire [95:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.TinyRocketConfig.fir 200785:4]
  wire [95:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.TinyRocketConfig.fir 200786:4]
  wire [383:0] a_opcodes_set = _GEN_19[383:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200570:4]
  wire [383:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.TinyRocketConfig.fir 200788:4]
  wire [383:0] d_opcodes_clr = _GEN_23[383:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200657:4]
  wire [383:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.TinyRocketConfig.fir 200789:4]
  wire [383:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.TinyRocketConfig.fir 200790:4]
  wire [383:0] a_sizes_set = _GEN_20[383:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200572:4]
  wire [383:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.TinyRocketConfig.fir 200792:4]
  wire [383:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.TinyRocketConfig.fir 200794:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 200796:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.TinyRocketConfig.fir 200799:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.TinyRocketConfig.fir 200800:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.TinyRocketConfig.fir 200801:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.TinyRocketConfig.fir 200802:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.TinyRocketConfig.fir 200803:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.TinyRocketConfig.fir 200804:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200806:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200807:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.TinyRocketConfig.fir 200813:4]
  wire  _T_676 = a_first_done | d_first_done; // @[Monitor.scala 712:27 chipyard.TestHarness.TinyRocketConfig.fir 200817:4]
  reg [95:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.TinyRocketConfig.fir 200821:4]
  reg [383:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 200823:4]
  reg  d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200858:4]
  wire  d_first_counter1_2 = d_first_counter_2 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 200860:4]
  wire  d_first_2 = ~d_first_counter_2; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 200861:4]
  wire [383:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.TinyRocketConfig.fir 200894:4]
  wire [383:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.TinyRocketConfig.fir 200899:4]
  wire [383:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[383:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.TinyRocketConfig.fir 200900:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.TinyRocketConfig.fir 200978:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.TinyRocketConfig.fir 200980:4]
  wire  _T_698 = d_first_done & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.TinyRocketConfig.fir 200986:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.TinyRocketConfig.fir 200988:4]
  wire [127:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.TinyRocketConfig.fir 200989:4 Monitor.scala 784:21 chipyard.TestHarness.TinyRocketConfig.fir 200991:6 chipyard.TestHarness.TinyRocketConfig.fir 200970:4]
  wire [1038:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.TinyRocketConfig.fir 200989:4 Monitor.scala 785:21 chipyard.TestHarness.TinyRocketConfig.fir 200998:6 chipyard.TestHarness.TinyRocketConfig.fir 200974:4]
  wire [95:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.TinyRocketConfig.fir 201024:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 201028:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 201029:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200882:4 Monitor.scala 747:21 chipyard.TestHarness.TinyRocketConfig.fir 200901:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.TinyRocketConfig.fir 201047:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 201049:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 201050:8]
  wire [95:0] d_clr_1 = _GEN_67[95:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200969:4]
  wire [95:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.TinyRocketConfig.fir 201092:4]
  wire [95:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.TinyRocketConfig.fir 201093:4]
  wire [383:0] d_opcodes_clr_1 = _GEN_68[383:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 200973:4]
  wire [383:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.TinyRocketConfig.fir 201096:4]
  wire [383:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.TinyRocketConfig.fir 201101:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.TinyRocketConfig.fir 201103:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.TinyRocketConfig.fir 201106:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.TinyRocketConfig.fir 201107:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.TinyRocketConfig.fir 201108:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.TinyRocketConfig.fir 201109:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.TinyRocketConfig.fir 201110:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.TinyRocketConfig.fir 201111:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 201113:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 201114:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.TinyRocketConfig.fir 201120:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199448:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199546:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199643:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199734:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199799:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199863:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199925:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199987:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200057:10]
  wire  _GEN_202 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200099:10]
  wire  _GEN_208 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200157:10]
  wire  _GEN_214 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200216:10]
  wire  _GEN_216 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200251:10]
  wire  _GEN_218 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200287:10]
  wire  _GEN_220 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200720:10]
  wire  _GEN_225 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200742:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 200797:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 201104:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200356:4]
      a_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200356:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 200366:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 200367:6]
        a_first_counter <= 1'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 200421:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.TinyRocketConfig.fir 200422:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 200421:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.TinyRocketConfig.fir 200423:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 200421:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.TinyRocketConfig.fir 200424:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 200421:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.TinyRocketConfig.fir 200425:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 200421:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.TinyRocketConfig.fir 200426:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200436:4]
      d_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200436:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 200446:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 200447:6]
        d_first_counter <= 1'h0;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 200510:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.TinyRocketConfig.fir 200511:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 200510:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.TinyRocketConfig.fir 200513:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 200510:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.TinyRocketConfig.fir 200514:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 200518:4]
      inflight <= 96'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 200518:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.TinyRocketConfig.fir 200787:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 200519:4]
      inflight_opcodes <= 384'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 200519:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.TinyRocketConfig.fir 200791:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 200520:4]
      inflight_sizes <= 384'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 200520:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.TinyRocketConfig.fir 200795:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200530:4]
      a_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200530:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 200540:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 200541:6]
        a_first_counter_1 <= 1'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200552:4]
      d_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200552:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 200562:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 200563:6]
        d_first_counter_1 <= 1'h0;
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 200796:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 200796:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.TinyRocketConfig.fir 200818:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.TinyRocketConfig.fir 200819:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.TinyRocketConfig.fir 200814:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.TinyRocketConfig.fir 200821:4]
      inflight_1 <= 96'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.TinyRocketConfig.fir 200821:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.TinyRocketConfig.fir 201094:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 200823:4]
      inflight_sizes_1 <= 384'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 200823:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.TinyRocketConfig.fir 201102:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200858:4]
      d_first_counter_2 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 200858:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 200868:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 200869:6]
        d_first_counter_2 <= 1'h0;
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.TinyRocketConfig.fir 201103:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.TinyRocketConfig.fir 201103:4]
    end else if (d_first_done) begin // @[Monitor.scala 819:47 chipyard.TestHarness.TinyRocketConfig.fir 201127:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.TinyRocketConfig.fir 201128:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.TinyRocketConfig.fir 201121:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199448:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199449:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199467:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199468:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199474:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199475:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199482:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199483:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199489:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199490:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199497:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199498:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199506:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199507:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199514:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199515:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199546:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199547:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199565:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199566:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199572:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199573:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199580:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199581:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199587:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199588:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199595:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199596:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199603:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199604:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199612:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199613:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199620:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199621:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199643:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199644:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199661:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199662:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199668:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199669:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199675:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199676:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199683:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199684:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199691:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199692:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199699:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199700:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199734:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199735:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199741:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199742:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199748:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199749:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199756:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199757:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199764:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199765:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199799:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199800:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199806:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199807:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199813:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199814:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199821:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199822:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199831:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199832:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199863:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199864:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199870:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199871:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199877:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199878:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199885:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199886:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199893:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199894:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199925:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199926:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199932:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199933:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199939:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199940:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199947:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199948:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199955:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199956:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199987:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199988:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199994:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 199995:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200001:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200002:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200009:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200010:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200017:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200018:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200025:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200026:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200036:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200037:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200057:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200058:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200065:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200066:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200099:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200100:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200106:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200107:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200114:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200115:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200157:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200158:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200164:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200165:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200172:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200173:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200216:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_214 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200217:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200251:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_216 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200252:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200287:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_218 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200288:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200383:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200384:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200391:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200392:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200399:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200400:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200407:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200408:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200415:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200416:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200464:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200465:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200480:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200481:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200488:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200489:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200649:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200650:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200709:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200710:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200720:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200721:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_220 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200728:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200729:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200742:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200743:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200750:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200751:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200769:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200770:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200781:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 200782:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200809:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 200810:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 201031:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 201032:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 201052:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 201053:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 201116:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 201117:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[6:0];
  _RAND_10 = {3{`RANDOM}};
  inflight = _RAND_10[95:0];
  _RAND_11 = {12{`RANDOM}};
  inflight_opcodes = _RAND_11[383:0];
  _RAND_12 = {12{`RANDOM}};
  inflight_sizes = _RAND_12[383:0];
  _RAND_13 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  watchdog = _RAND_15[31:0];
  _RAND_16 = {3{`RANDOM}};
  inflight_1 = _RAND_16[95:0];
  _RAND_17 = {12{`RANDOM}};
  inflight_sizes_1 = _RAND_17[383:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  watchdog_1 = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLRAM_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 201131:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 201132:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 201133:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  input  [1:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  input  [6:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  input  [3:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  input  [31:0] auto_in_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  output [1:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  output [6:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
  output [31:0] auto_in_d_bits_data // @[chipyard.TestHarness.TinyRocketConfig.fir 201134:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire [1:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire [6:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire [1:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire [6:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
  wire [9:0] mem_RW0_addr; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire  mem_RW0_en; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire  mem_RW0_clk; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire  mem_RW0_wmode; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire [7:0] mem_RW0_wdata_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire [7:0] mem_RW0_wdata_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire [7:0] mem_RW0_wdata_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire [7:0] mem_RW0_wdata_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire [7:0] mem_RW0_rdata_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire [7:0] mem_RW0_rdata_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire [7:0] mem_RW0_rdata_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire [7:0] mem_RW0_rdata_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire  mem_RW0_wmask_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire  mem_RW0_wmask_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire  mem_RW0_wmask_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  wire  mem_RW0_wmask_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
  reg  r_full; // @[SRAM.scala 134:30 chipyard.TestHarness.TinyRocketConfig.fir 201180:4]
  reg [1:0] r_size; // @[SRAM.scala 137:26 chipyard.TestHarness.TinyRocketConfig.fir 201183:4]
  reg [6:0] r_source; // @[SRAM.scala 138:26 chipyard.TestHarness.TinyRocketConfig.fir 201184:4]
  reg  r_read; // @[SRAM.scala 139:26 chipyard.TestHarness.TinyRocketConfig.fir 201185:4]
  reg  REG; // @[SRAM.scala 321:58 chipyard.TestHarness.TinyRocketConfig.fir 201547:4]
  reg [7:0] r_1; // @[Reg.scala 15:16 chipyard.TestHarness.TinyRocketConfig.fir 201549:4]
  wire [7:0] r_raw_data_1 = REG ? mem_RW0_rdata_1 : r_1; // @[package.scala 79:42 chipyard.TestHarness.TinyRocketConfig.fir 201556:4]
  reg [7:0] r_0; // @[Reg.scala 15:16 chipyard.TestHarness.TinyRocketConfig.fir 201549:4]
  wire [7:0] r_raw_data_0 = REG ? mem_RW0_rdata_0 : r_0; // @[package.scala 79:42 chipyard.TestHarness.TinyRocketConfig.fir 201556:4]
  wire [15:0] r_corrected_lo = {r_raw_data_1,r_raw_data_0}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 201218:4]
  reg [7:0] r_3; // @[Reg.scala 15:16 chipyard.TestHarness.TinyRocketConfig.fir 201549:4]
  wire [7:0] r_raw_data_3 = REG ? mem_RW0_rdata_3 : r_3; // @[package.scala 79:42 chipyard.TestHarness.TinyRocketConfig.fir 201556:4]
  reg [7:0] r_2; // @[Reg.scala 15:16 chipyard.TestHarness.TinyRocketConfig.fir 201549:4]
  wire [7:0] r_raw_data_2 = REG ? mem_RW0_rdata_2 : r_2; // @[package.scala 79:42 chipyard.TestHarness.TinyRocketConfig.fir 201556:4]
  wire [15:0] r_corrected_hi = {r_raw_data_3,r_raw_data_2}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 201219:4]
  wire  _bundleIn_0_a_ready_T_2 = ~r_full; // @[SRAM.scala 243:41 chipyard.TestHarness.TinyRocketConfig.fir 201347:4]
  wire  in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.TinyRocketConfig.fir 201348:4]
  wire  a_read = auto_in_a_bits_opcode == 3'h4; // @[SRAM.scala 251:35 chipyard.TestHarness.TinyRocketConfig.fir 201356:4]
  wire  _GEN_18 = auto_in_d_ready ? 1'h0 : r_full; // @[SRAM.scala 273:20 chipyard.TestHarness.TinyRocketConfig.fir 201381:4 SRAM.scala 273:29 chipyard.TestHarness.TinyRocketConfig.fir 201382:6 SRAM.scala 134:30 chipyard.TestHarness.TinyRocketConfig.fir 201180:4]
  wire  _T_18 = in_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 201384:4]
  wire  _T_19 = ~a_read; // @[SRAM.scala 287:13 chipyard.TestHarness.TinyRocketConfig.fir 201398:6]
  wire  _GEN_20 = _T_18 | _GEN_18; // @[SRAM.scala 274:24 chipyard.TestHarness.TinyRocketConfig.fir 201385:4 SRAM.scala 275:18 chipyard.TestHarness.TinyRocketConfig.fir 201386:6]
  wire  a_lanes_lo_lo = |auto_in_a_bits_mask[0]; // @[SRAM.scala 303:95 chipyard.TestHarness.TinyRocketConfig.fir 201466:4]
  wire  a_lanes_lo_hi = |auto_in_a_bits_mask[1]; // @[SRAM.scala 303:95 chipyard.TestHarness.TinyRocketConfig.fir 201468:4]
  wire  a_lanes_hi_lo = |auto_in_a_bits_mask[2]; // @[SRAM.scala 303:95 chipyard.TestHarness.TinyRocketConfig.fir 201470:4]
  wire  a_lanes_hi_hi = |auto_in_a_bits_mask[3]; // @[SRAM.scala 303:95 chipyard.TestHarness.TinyRocketConfig.fir 201472:4]
  wire [3:0] a_lanes = {a_lanes_hi_hi,a_lanes_hi_lo,a_lanes_lo_hi,a_lanes_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 201475:4]
  wire  wen = _T_18 & _T_19; // @[SRAM.scala 309:52 chipyard.TestHarness.TinyRocketConfig.fir 201483:4]
  wire  _ren_T = ~wen; // @[SRAM.scala 310:15 chipyard.TestHarness.TinyRocketConfig.fir 201486:4]
  wire  ren = _ren_T & _T_18; // @[SRAM.scala 310:20 chipyard.TestHarness.TinyRocketConfig.fir 201488:4]
  wire  index_lo_lo_lo = auto_in_a_bits_address[2]; // @[SRAM.scala 320:60 chipyard.TestHarness.TinyRocketConfig.fir 201503:4]
  wire  index_lo_lo_hi = auto_in_a_bits_address[3]; // @[SRAM.scala 320:60 chipyard.TestHarness.TinyRocketConfig.fir 201504:4]
  wire  index_lo_hi_lo = auto_in_a_bits_address[4]; // @[SRAM.scala 320:60 chipyard.TestHarness.TinyRocketConfig.fir 201505:4]
  wire  index_lo_hi_hi_lo = auto_in_a_bits_address[5]; // @[SRAM.scala 320:60 chipyard.TestHarness.TinyRocketConfig.fir 201506:4]
  wire  index_lo_hi_hi_hi = auto_in_a_bits_address[6]; // @[SRAM.scala 320:60 chipyard.TestHarness.TinyRocketConfig.fir 201507:4]
  wire  index_hi_lo_lo = auto_in_a_bits_address[7]; // @[SRAM.scala 320:60 chipyard.TestHarness.TinyRocketConfig.fir 201508:4]
  wire  index_hi_lo_hi = auto_in_a_bits_address[8]; // @[SRAM.scala 320:60 chipyard.TestHarness.TinyRocketConfig.fir 201509:4]
  wire  index_hi_hi_lo = auto_in_a_bits_address[9]; // @[SRAM.scala 320:60 chipyard.TestHarness.TinyRocketConfig.fir 201510:4]
  wire  index_hi_hi_hi_lo = auto_in_a_bits_address[10]; // @[SRAM.scala 320:60 chipyard.TestHarness.TinyRocketConfig.fir 201511:4]
  wire  index_hi_hi_hi_hi = auto_in_a_bits_address[11]; // @[SRAM.scala 320:60 chipyard.TestHarness.TinyRocketConfig.fir 201512:4]
  wire [4:0] index_lo = {index_lo_hi_hi_hi,index_lo_hi_hi_lo,index_lo_hi_lo,index_lo_lo_hi,index_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 201533:4]
  wire [4:0] index_hi = {index_hi_hi_hi_hi,index_hi_hi_hi_lo,index_hi_hi_lo,index_hi_lo_hi,index_hi_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 201537:4]
  TLMonitor_42_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 201141:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source)
  );
  mem_inTestHarness mem ( // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.TinyRocketConfig.fir 201165:4]
    .RW0_addr(mem_RW0_addr),
    .RW0_en(mem_RW0_en),
    .RW0_clk(mem_RW0_clk),
    .RW0_wmode(mem_RW0_wmode),
    .RW0_wdata_0(mem_RW0_wdata_0),
    .RW0_wdata_1(mem_RW0_wdata_1),
    .RW0_wdata_2(mem_RW0_wdata_2),
    .RW0_wdata_3(mem_RW0_wdata_3),
    .RW0_rdata_0(mem_RW0_rdata_0),
    .RW0_rdata_1(mem_RW0_rdata_1),
    .RW0_rdata_2(mem_RW0_rdata_2),
    .RW0_rdata_3(mem_RW0_rdata_3),
    .RW0_wmask_0(mem_RW0_wmask_0),
    .RW0_wmask_1(mem_RW0_wmask_1),
    .RW0_wmask_2(mem_RW0_wmask_2),
    .RW0_wmask_3(mem_RW0_wmask_3)
  );
  assign auto_in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.TinyRocketConfig.fir 201348:4]
  assign auto_in_d_valid = r_full; // @[SRAM.scala 240:65 chipyard.TestHarness.TinyRocketConfig.fir 201327:4]
  assign auto_in_d_bits_opcode = {{2'd0}, r_read}; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 SRAM.scala 209:23 chipyard.TestHarness.TinyRocketConfig.fir 201275:4]
  assign auto_in_d_bits_size = r_size; // @[SRAM.scala 211:29 chipyard.TestHarness.TinyRocketConfig.fir 201277:4]
  assign auto_in_d_bits_source = r_source; // @[SRAM.scala 212:29 chipyard.TestHarness.TinyRocketConfig.fir 201279:4]
  assign auto_in_d_bits_data = {r_corrected_hi,r_corrected_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 201223:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 201142:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 201143:4]
  assign monitor_io_in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.TinyRocketConfig.fir 201348:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201164:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201164:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201164:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201164:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201164:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201164:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201164:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201164:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201164:4]
  assign monitor_io_in_d_valid = r_full; // @[SRAM.scala 240:65 chipyard.TestHarness.TinyRocketConfig.fir 201327:4]
  assign monitor_io_in_d_bits_opcode = {{2'd0}, r_read}; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201139:4 SRAM.scala 209:23 chipyard.TestHarness.TinyRocketConfig.fir 201275:4]
  assign monitor_io_in_d_bits_size = r_size; // @[SRAM.scala 211:29 chipyard.TestHarness.TinyRocketConfig.fir 201277:4]
  assign monitor_io_in_d_bits_source = r_source; // @[SRAM.scala 212:29 chipyard.TestHarness.TinyRocketConfig.fir 201279:4]
  assign mem_RW0_wdata_0 = auto_in_a_bits_data[7:0]; // @[SRAM.scala 291:67 chipyard.TestHarness.TinyRocketConfig.fir 201403:4]
  assign mem_RW0_wdata_1 = auto_in_a_bits_data[15:8]; // @[SRAM.scala 291:67 chipyard.TestHarness.TinyRocketConfig.fir 201404:4]
  assign mem_RW0_wdata_2 = auto_in_a_bits_data[23:16]; // @[SRAM.scala 291:67 chipyard.TestHarness.TinyRocketConfig.fir 201405:4]
  assign mem_RW0_wdata_3 = auto_in_a_bits_data[31:24]; // @[SRAM.scala 291:67 chipyard.TestHarness.TinyRocketConfig.fir 201406:4]
  assign mem_RW0_wmask_0 = a_lanes[0]; // @[SRAM.scala 322:46 chipyard.TestHarness.TinyRocketConfig.fir 201562:6]
  assign mem_RW0_wmask_1 = a_lanes[1]; // @[SRAM.scala 322:46 chipyard.TestHarness.TinyRocketConfig.fir 201563:6]
  assign mem_RW0_wmask_2 = a_lanes[2]; // @[SRAM.scala 322:46 chipyard.TestHarness.TinyRocketConfig.fir 201564:6]
  assign mem_RW0_wmask_3 = a_lanes[3]; // @[SRAM.scala 322:46 chipyard.TestHarness.TinyRocketConfig.fir 201565:6]
  assign mem_RW0_wmode = _T_18 & _T_19; // @[SRAM.scala 309:52 chipyard.TestHarness.TinyRocketConfig.fir 201483:4]
  assign mem_RW0_clk = clock;
  assign mem_RW0_en = ren | wen;
  assign mem_RW0_addr = {index_hi,index_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 201538:4]
  always @(posedge clock) begin
    if (reset) begin // @[SRAM.scala 134:30 chipyard.TestHarness.TinyRocketConfig.fir 201180:4]
      r_full <= 1'h0; // @[SRAM.scala 134:30 chipyard.TestHarness.TinyRocketConfig.fir 201180:4]
    end else begin
      r_full <= _GEN_20;
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.TinyRocketConfig.fir 201385:4]
      r_size <= auto_in_a_bits_size; // @[SRAM.scala 279:18 chipyard.TestHarness.TinyRocketConfig.fir 201390:6]
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.TinyRocketConfig.fir 201385:4]
      r_source <= auto_in_a_bits_source; // @[SRAM.scala 280:18 chipyard.TestHarness.TinyRocketConfig.fir 201391:6]
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.TinyRocketConfig.fir 201385:4]
      r_read <= a_read; // @[SRAM.scala 281:18 chipyard.TestHarness.TinyRocketConfig.fir 201392:6]
    end
    REG <= _ren_T & _T_18; // @[SRAM.scala 310:20 chipyard.TestHarness.TinyRocketConfig.fir 201488:4]
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.TinyRocketConfig.fir 201550:4]
      r_1 <= mem_RW0_rdata_1; // @[Reg.scala 16:23 chipyard.TestHarness.TinyRocketConfig.fir 201552:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.TinyRocketConfig.fir 201550:4]
      r_0 <= mem_RW0_rdata_0; // @[Reg.scala 16:23 chipyard.TestHarness.TinyRocketConfig.fir 201551:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.TinyRocketConfig.fir 201550:4]
      r_3 <= mem_RW0_rdata_3; // @[Reg.scala 16:23 chipyard.TestHarness.TinyRocketConfig.fir 201554:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.TinyRocketConfig.fir 201550:4]
      r_2 <= mem_RW0_rdata_2; // @[Reg.scala 16:23 chipyard.TestHarness.TinyRocketConfig.fir 201553:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_size = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  r_source = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  r_read = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  r_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  r_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  r_2 = _RAND_8[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar_9_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 201590:2]
  output        auto_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [2:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [1:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [3:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [31:0] auto_in_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [2:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [1:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [31:0] auto_in_d_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [2:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [1:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [3:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output [31:0] auto_out_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [2:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [1:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input         auto_out_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input  [31:0] auto_out_d_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 201593:4]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 201598:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 201602:4]
  assign auto_in_d_valid = auto_out_d_valid; // @[ReadyValidCancel.scala 21:38 chipyard.TestHarness.TinyRocketConfig.fir 202014:4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 201598:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 201602:4]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 201598:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 201602:4]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 201598:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 201602:4]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Xbar.scala 228:69 chipyard.TestHarness.TinyRocketConfig.fir 201713:4]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Xbar.scala 323:53 chipyard.TestHarness.TinyRocketConfig.fir 201775:4]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 201598:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 201602:4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 201598:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 201602:4]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 201598:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 201602:4]
  assign auto_out_a_valid = auto_in_a_valid; // @[ReadyValidCancel.scala 21:38 chipyard.TestHarness.TinyRocketConfig.fir 202039:4]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201600:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201603:4]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201600:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201603:4]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201600:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201603:4]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55 chipyard.TestHarness.TinyRocketConfig.fir 201667:4]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201600:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201603:4]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201600:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201603:4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201600:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201603:4]
  assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201600:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201603:4]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 201600:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 201603:4]
endmodule
module TLMonitor_43_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 202116:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 202117:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 202118:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input  [1:0]  io_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input  [6:0]  io_in_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input  [3:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input  [1:0]  io_in_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input  [6:0]  io_in_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input         io_in_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 202119:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [95:0] _RAND_13;
  reg [383:0] _RAND_14;
  reg [383:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [95:0] _RAND_19;
  reg [383:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 203579:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 203886:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 7'h5f; // @[Parameters.scala 57:20 chipyard.TestHarness.TinyRocketConfig.fir 202136:6]
  wire [4:0] _is_aligned_mask_T_1 = 5'h3 << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 202142:6]
  wire [1:0] is_aligned_mask = ~_is_aligned_mask_T_1[1:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 202144:6]
  wire [28:0] _GEN_71 = {{27'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.TinyRocketConfig.fir 202145:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.TinyRocketConfig.fir 202145:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.TinyRocketConfig.fir 202146:6]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49 chipyard.TestHarness.TinyRocketConfig.fir 202148:6]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.TinyRocketConfig.fir 202149:6]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81 chipyard.TestHarness.TinyRocketConfig.fir 202151:6]
  wire  _mask_T = io_in_a_bits_size >= 2'h2; // @[Misc.scala 205:21 chipyard.TestHarness.TinyRocketConfig.fir 202152:6]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 202153:6]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 202154:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 202155:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 202157:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 202158:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 202160:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 202161:6]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 202162:6]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 202163:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 202164:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 202165:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 202166:6]
  wire  mask_lo_lo = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 202167:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 202168:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 202169:6]
  wire  mask_lo_hi = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 202170:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 202171:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 202172:6]
  wire  mask_hi_lo = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 202173:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 202174:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 202175:6]
  wire  mask_hi_hi = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 202176:6]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 202179:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.TinyRocketConfig.fir 202202:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 202218:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 202219:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 202221:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 202222:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202228:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202253:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202254:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202261:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202262:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202268:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202269:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.TinyRocketConfig.fir 202274:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202276:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202277:8]
  wire [3:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.TinyRocketConfig.fir 202282:8]
  wire  _T_74 = _T_73 == 4'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.TinyRocketConfig.fir 202283:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202285:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202286:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.TinyRocketConfig.fir 202291:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202293:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202294:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.TinyRocketConfig.fir 202300:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.TinyRocketConfig.fir 202380:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202382:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202383:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.TinyRocketConfig.fir 202406:6]
  wire  _T_164 = io_in_a_bits_size <= 2'h2; // @[Parameters.scala 92:42 chipyard.TestHarness.TinyRocketConfig.fir 202429:8]
  wire  _T_172 = _T_164 & _T_37; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 202437:8]
  wire  _T_175 = _T_172 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202440:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202441:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.TinyRocketConfig.fir 202460:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202462:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202463:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.TinyRocketConfig.fir 202468:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202470:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202471:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.TinyRocketConfig.fir 202485:6]
  wire  _T_218 = _source_ok_T_4 & _T_172; // @[Monitor.scala 115:71 chipyard.TestHarness.TinyRocketConfig.fir 202511:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202513:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202514:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.TinyRocketConfig.fir 202550:6]
  wire [3:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.TinyRocketConfig.fir 202606:8]
  wire [3:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.TinyRocketConfig.fir 202607:8]
  wire  _T_275 = _T_274 == 4'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.TinyRocketConfig.fir 202608:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202610:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202611:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.TinyRocketConfig.fir 202617:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.TinyRocketConfig.fir 202662:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202664:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202665:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.TinyRocketConfig.fir 202679:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.TinyRocketConfig.fir 202724:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202726:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202727:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.TinyRocketConfig.fir 202741:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.TinyRocketConfig.fir 202786:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202788:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202789:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.TinyRocketConfig.fir 202813:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202815:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202816:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 7'h5f; // @[Parameters.scala 57:20 chipyard.TestHarness.TinyRocketConfig.fir 202827:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.TinyRocketConfig.fir 202833:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202836:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202837:8]
  wire  _T_405 = io_in_d_bits_size >= 2'h2; // @[Monitor.scala 312:27 chipyard.TestHarness.TinyRocketConfig.fir 202842:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202844:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202845:8]
  wire  _T_409 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.TinyRocketConfig.fir 202850:8]
  wire  _T_411 = _T_409 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202852:8]
  wire  _T_412 = ~_T_411; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202853:8]
  wire  _T_413 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.TinyRocketConfig.fir 202858:8]
  wire  _T_415 = _T_413 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202860:8]
  wire  _T_416 = ~_T_415; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202861:8]
  wire  _T_417 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.TinyRocketConfig.fir 202866:8]
  wire  _T_419 = _T_417 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202868:8]
  wire  _T_420 = ~_T_419; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202869:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.TinyRocketConfig.fir 202875:6]
  wire  _T_432 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.TinyRocketConfig.fir 202899:8]
  wire  _T_434 = _T_432 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202901:8]
  wire  _T_435 = ~_T_434; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202902:8]
  wire  _T_436 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.TinyRocketConfig.fir 202907:8]
  wire  _T_438 = _T_436 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202909:8]
  wire  _T_439 = ~_T_438; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202910:8]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.TinyRocketConfig.fir 202933:6]
  wire  _T_469 = _T_417 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.TinyRocketConfig.fir 202974:8]
  wire  _T_471 = _T_469 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202976:8]
  wire  _T_472 = ~_T_471; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202977:8]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.TinyRocketConfig.fir 202992:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.TinyRocketConfig.fir 203027:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.TinyRocketConfig.fir 203063:6]
  wire  a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 203129:4]
  reg  a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203138:4]
  wire  a_first_counter1 = a_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 203140:4]
  wire  a_first = ~a_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 203141:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.TinyRocketConfig.fir 203152:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.TinyRocketConfig.fir 203153:4]
  reg [1:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.TinyRocketConfig.fir 203154:4]
  reg [6:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.TinyRocketConfig.fir 203155:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.TinyRocketConfig.fir 203156:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.TinyRocketConfig.fir 203157:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.TinyRocketConfig.fir 203158:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.TinyRocketConfig.fir 203160:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203162:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203163:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.TinyRocketConfig.fir 203168:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203170:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203171:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.TinyRocketConfig.fir 203176:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203178:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203179:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.TinyRocketConfig.fir 203184:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203186:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203187:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.TinyRocketConfig.fir 203192:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203194:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203195:6]
  wire  _T_565 = a_first_done & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.TinyRocketConfig.fir 203202:4]
  wire  d_first_done = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 203210:4]
  reg  d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203218:4]
  wire  d_first_counter1 = d_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 203220:4]
  wire  d_first = ~d_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 203221:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.TinyRocketConfig.fir 203232:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.TinyRocketConfig.fir 203233:4]
  reg [1:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.TinyRocketConfig.fir 203234:4]
  reg [6:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.TinyRocketConfig.fir 203235:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.TinyRocketConfig.fir 203236:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.TinyRocketConfig.fir 203237:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.TinyRocketConfig.fir 203238:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.TinyRocketConfig.fir 203239:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.TinyRocketConfig.fir 203241:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203243:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203244:6]
  wire  _T_572 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.TinyRocketConfig.fir 203249:6]
  wire  _T_574 = _T_572 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203251:6]
  wire  _T_575 = ~_T_574; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203252:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.TinyRocketConfig.fir 203257:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203259:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203260:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.TinyRocketConfig.fir 203265:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203267:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203268:6]
  wire  _T_584 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.TinyRocketConfig.fir 203273:6]
  wire  _T_586 = _T_584 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203275:6]
  wire  _T_587 = ~_T_586; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203276:6]
  wire  _T_588 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.TinyRocketConfig.fir 203281:6]
  wire  _T_590 = _T_588 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203283:6]
  wire  _T_591 = ~_T_590; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203284:6]
  wire  _T_593 = d_first_done & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.TinyRocketConfig.fir 203291:4]
  reg [95:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 203300:4]
  reg [383:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 203301:4]
  reg [383:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 203302:4]
  reg  a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203312:4]
  wire  a_first_counter1_1 = a_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 203314:4]
  wire  a_first_1 = ~a_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 203315:4]
  reg  d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203334:4]
  wire  d_first_counter1_1 = d_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 203336:4]
  wire  d_first_1 = ~d_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 203337:4]
  wire [8:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.TinyRocketConfig.fir 203358:4]
  wire [9:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.TinyRocketConfig.fir 203358:4]
  wire [383:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.TinyRocketConfig.fir 203359:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.TinyRocketConfig.fir 203363:4]
  wire [383:0] _GEN_73 = {{368'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.TinyRocketConfig.fir 203364:4]
  wire [383:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.TinyRocketConfig.fir 203364:4]
  wire [383:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[383:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.TinyRocketConfig.fir 203365:4]
  wire [383:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.TinyRocketConfig.fir 203370:4]
  wire [383:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.TinyRocketConfig.fir 203375:4]
  wire [383:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[383:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.TinyRocketConfig.fir 203376:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.TinyRocketConfig.fir 203400:4]
  wire [127:0] _a_set_wo_ready_T = 128'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.TinyRocketConfig.fir 203403:6]
  wire [127:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.TinyRocketConfig.fir 203402:4 Monitor.scala 649:22 chipyard.TestHarness.TinyRocketConfig.fir 203404:6 chipyard.TestHarness.TinyRocketConfig.fir 203351:4]
  wire  _T_597 = a_first_done & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.TinyRocketConfig.fir 203407:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.TinyRocketConfig.fir 203412:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.TinyRocketConfig.fir 203413:6]
  wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.TinyRocketConfig.fir 203415:6]
  wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.TinyRocketConfig.fir 203416:6]
  wire [8:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.TinyRocketConfig.fir 203418:6]
  wire [9:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.TinyRocketConfig.fir 203418:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 203409:4 Monitor.scala 654:28 chipyard.TestHarness.TinyRocketConfig.fir 203414:6 chipyard.TestHarness.TinyRocketConfig.fir 203397:4]
  wire [1026:0] _GEN_79 = {{1023'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.TinyRocketConfig.fir 203419:6]
  wire [1026:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.TinyRocketConfig.fir 203419:6]
  wire [2:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 3'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 203409:4 Monitor.scala 655:28 chipyard.TestHarness.TinyRocketConfig.fir 203417:6 chipyard.TestHarness.TinyRocketConfig.fir 203399:4]
  wire [1025:0] _GEN_81 = {{1023'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.TinyRocketConfig.fir 203422:6]
  wire [1025:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.TinyRocketConfig.fir 203422:6]
  wire [95:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.TinyRocketConfig.fir 203424:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.TinyRocketConfig.fir 203426:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203428:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203429:6]
  wire [127:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 128'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 203409:4 Monitor.scala 653:28 chipyard.TestHarness.TinyRocketConfig.fir 203411:6 chipyard.TestHarness.TinyRocketConfig.fir 203349:4]
  wire [1026:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 1027'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 203409:4 Monitor.scala 656:28 chipyard.TestHarness.TinyRocketConfig.fir 203420:6 chipyard.TestHarness.TinyRocketConfig.fir 203353:4]
  wire [1025:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 1026'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 203409:4 Monitor.scala 657:28 chipyard.TestHarness.TinyRocketConfig.fir 203423:6 chipyard.TestHarness.TinyRocketConfig.fir 203355:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.TinyRocketConfig.fir 203444:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.TinyRocketConfig.fir 203446:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.TinyRocketConfig.fir 203447:4]
  wire [127:0] _d_clr_wo_ready_T = 128'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.TinyRocketConfig.fir 203449:6]
  wire [127:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.TinyRocketConfig.fir 203448:4 Monitor.scala 672:22 chipyard.TestHarness.TinyRocketConfig.fir 203450:6 chipyard.TestHarness.TinyRocketConfig.fir 203438:4]
  wire  _T_610 = d_first_done & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.TinyRocketConfig.fir 203453:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.TinyRocketConfig.fir 203456:4]
  wire [1038:0] _GEN_83 = {{1023'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.TinyRocketConfig.fir 203465:6]
  wire [1038:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.TinyRocketConfig.fir 203465:6]
  wire [127:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 203457:4 Monitor.scala 676:21 chipyard.TestHarness.TinyRocketConfig.fir 203459:6 chipyard.TestHarness.TinyRocketConfig.fir 203436:4]
  wire [1038:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 203457:4 Monitor.scala 677:21 chipyard.TestHarness.TinyRocketConfig.fir 203466:6 chipyard.TestHarness.TinyRocketConfig.fir 203440:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.TinyRocketConfig.fir 203482:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.TinyRocketConfig.fir 203483:6]
  wire [95:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.TinyRocketConfig.fir 203484:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.TinyRocketConfig.fir 203486:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203488:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203489:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 203495:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 203496:8 Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 203496:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 203496:8 Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 203496:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 203496:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.TinyRocketConfig.fir 203497:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203499:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203500:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.TinyRocketConfig.fir 203505:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203507:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203508:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203356:4 Monitor.scala 634:21 chipyard.TestHarness.TinyRocketConfig.fir 203366:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 203516:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 203518:8 Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 203518:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 203518:8 Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 203518:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 203518:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.TinyRocketConfig.fir 203519:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203521:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203522:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203367:4 Monitor.scala 638:19 chipyard.TestHarness.TinyRocketConfig.fir 203377:4]
  wire [3:0] _GEN_86 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.TinyRocketConfig.fir 203527:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.TinyRocketConfig.fir 203527:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203529:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203530:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.TinyRocketConfig.fir 203538:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.TinyRocketConfig.fir 203539:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.TinyRocketConfig.fir 203541:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.TinyRocketConfig.fir 203543:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.TinyRocketConfig.fir 203545:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.TinyRocketConfig.fir 203546:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203548:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203549:6]
  wire [95:0] a_set_wo_ready = _GEN_15[95:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203350:4]
  wire [95:0] d_clr_wo_ready = _GEN_21[95:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203437:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.TinyRocketConfig.fir 203555:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.TinyRocketConfig.fir 203556:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.TinyRocketConfig.fir 203557:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.TinyRocketConfig.fir 203558:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203560:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203561:4]
  wire [95:0] a_set = _GEN_16[95:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203348:4]
  wire [95:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.TinyRocketConfig.fir 203566:4]
  wire [95:0] d_clr = _GEN_22[95:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203435:4]
  wire [95:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.TinyRocketConfig.fir 203567:4]
  wire [95:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.TinyRocketConfig.fir 203568:4]
  wire [383:0] a_opcodes_set = _GEN_19[383:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203352:4]
  wire [383:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.TinyRocketConfig.fir 203570:4]
  wire [383:0] d_opcodes_clr = _GEN_23[383:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203439:4]
  wire [383:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.TinyRocketConfig.fir 203571:4]
  wire [383:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.TinyRocketConfig.fir 203572:4]
  wire [383:0] a_sizes_set = _GEN_20[383:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203354:4]
  wire [383:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.TinyRocketConfig.fir 203574:4]
  wire [383:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.TinyRocketConfig.fir 203576:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 203578:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.TinyRocketConfig.fir 203581:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.TinyRocketConfig.fir 203582:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.TinyRocketConfig.fir 203583:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.TinyRocketConfig.fir 203584:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.TinyRocketConfig.fir 203585:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.TinyRocketConfig.fir 203586:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203588:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203589:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.TinyRocketConfig.fir 203595:4]
  wire  _T_676 = a_first_done | d_first_done; // @[Monitor.scala 712:27 chipyard.TestHarness.TinyRocketConfig.fir 203599:4]
  reg [95:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.TinyRocketConfig.fir 203603:4]
  reg [383:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 203605:4]
  reg  d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203640:4]
  wire  d_first_counter1_2 = d_first_counter_2 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 203642:4]
  wire  d_first_2 = ~d_first_counter_2; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 203643:4]
  wire [383:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.TinyRocketConfig.fir 203676:4]
  wire [383:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.TinyRocketConfig.fir 203681:4]
  wire [383:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[383:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.TinyRocketConfig.fir 203682:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.TinyRocketConfig.fir 203760:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.TinyRocketConfig.fir 203762:4]
  wire  _T_698 = d_first_done & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.TinyRocketConfig.fir 203768:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.TinyRocketConfig.fir 203770:4]
  wire [127:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 128'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.TinyRocketConfig.fir 203771:4 Monitor.scala 784:21 chipyard.TestHarness.TinyRocketConfig.fir 203773:6 chipyard.TestHarness.TinyRocketConfig.fir 203752:4]
  wire [1038:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 1039'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.TinyRocketConfig.fir 203771:4 Monitor.scala 785:21 chipyard.TestHarness.TinyRocketConfig.fir 203780:6 chipyard.TestHarness.TinyRocketConfig.fir 203756:4]
  wire [95:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.TinyRocketConfig.fir 203806:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203810:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203811:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203664:4 Monitor.scala 747:21 chipyard.TestHarness.TinyRocketConfig.fir 203683:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.TinyRocketConfig.fir 203829:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203831:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203832:8]
  wire [95:0] d_clr_1 = _GEN_67[95:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203751:4]
  wire [95:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.TinyRocketConfig.fir 203874:4]
  wire [95:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.TinyRocketConfig.fir 203875:4]
  wire [383:0] d_opcodes_clr_1 = _GEN_68[383:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 203755:4]
  wire [383:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.TinyRocketConfig.fir 203878:4]
  wire [383:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.TinyRocketConfig.fir 203883:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.TinyRocketConfig.fir 203885:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.TinyRocketConfig.fir 203888:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.TinyRocketConfig.fir 203889:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.TinyRocketConfig.fir 203890:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.TinyRocketConfig.fir 203891:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.TinyRocketConfig.fir 203892:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.TinyRocketConfig.fir 203893:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203895:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203896:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.TinyRocketConfig.fir 203902:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202230:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202328:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202425:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202516:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202581:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202645:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202707:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202769:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202839:10]
  wire  _GEN_208 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202881:10]
  wire  _GEN_222 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202939:10]
  wire  _GEN_236 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202998:10]
  wire  _GEN_244 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203033:10]
  wire  _GEN_252 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203069:10]
  wire  _GEN_260 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203502:10]
  wire  _GEN_265 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203524:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 203579:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 203886:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203138:4]
      a_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203138:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 203148:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 203149:6]
        a_first_counter <= 1'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 203203:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.TinyRocketConfig.fir 203204:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 203203:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.TinyRocketConfig.fir 203205:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 203203:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.TinyRocketConfig.fir 203206:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 203203:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.TinyRocketConfig.fir 203207:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 203203:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.TinyRocketConfig.fir 203208:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203218:4]
      d_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203218:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 203228:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 203229:6]
        d_first_counter <= 1'h0;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 203292:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.TinyRocketConfig.fir 203293:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 203292:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.TinyRocketConfig.fir 203294:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 203292:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.TinyRocketConfig.fir 203295:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 203292:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.TinyRocketConfig.fir 203296:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 203292:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.TinyRocketConfig.fir 203297:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 203292:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.TinyRocketConfig.fir 203298:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 203300:4]
      inflight <= 96'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 203300:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.TinyRocketConfig.fir 203569:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 203301:4]
      inflight_opcodes <= 384'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 203301:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.TinyRocketConfig.fir 203573:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 203302:4]
      inflight_sizes <= 384'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 203302:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.TinyRocketConfig.fir 203577:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203312:4]
      a_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203312:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 203322:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 203323:6]
        a_first_counter_1 <= 1'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203334:4]
      d_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203334:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 203344:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 203345:6]
        d_first_counter_1 <= 1'h0;
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 203578:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 203578:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.TinyRocketConfig.fir 203600:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.TinyRocketConfig.fir 203601:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.TinyRocketConfig.fir 203596:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.TinyRocketConfig.fir 203603:4]
      inflight_1 <= 96'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.TinyRocketConfig.fir 203603:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.TinyRocketConfig.fir 203876:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 203605:4]
      inflight_sizes_1 <= 384'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 203605:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.TinyRocketConfig.fir 203884:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203640:4]
      d_first_counter_2 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 203640:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 203650:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 203651:6]
        d_first_counter_2 <= 1'h0;
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.TinyRocketConfig.fir 203885:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.TinyRocketConfig.fir 203885:4]
    end else if (d_first_done) begin // @[Monitor.scala 819:47 chipyard.TestHarness.TinyRocketConfig.fir 203909:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.TinyRocketConfig.fir 203910:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.TinyRocketConfig.fir 203903:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202230:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202231:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202249:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202250:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202256:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202257:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202264:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202265:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202271:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202272:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202279:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202280:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202288:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202289:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202296:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202297:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202328:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202329:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202347:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202348:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202354:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202355:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202362:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202363:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202369:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202370:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202377:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202378:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202385:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202386:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202394:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202395:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202402:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202403:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202425:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202426:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202443:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202444:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202450:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202451:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202457:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202458:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202465:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202466:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202473:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202474:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202481:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202482:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202516:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202517:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202523:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202524:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202530:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202531:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202538:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202539:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202546:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202547:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202581:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202582:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202588:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202589:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202595:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202596:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202603:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202604:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202613:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202614:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202645:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202646:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202652:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202653:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202659:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202660:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202667:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202668:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202675:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202676:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202707:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202708:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202714:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202715:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202721:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202722:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202729:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202730:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202737:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202738:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202769:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202770:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202776:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202777:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202783:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202784:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202791:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202792:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202799:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202800:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202807:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 202808:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202818:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202819:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202839:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202840:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202847:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202848:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202855:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202856:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202863:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202864:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202871:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202872:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202881:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202882:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202888:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202889:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202896:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202897:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202904:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202905:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202912:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202913:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202920:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202921:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202929:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202930:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202939:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202940:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202946:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202947:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202954:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202955:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202962:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202963:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202970:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202971:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202979:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202980:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202988:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202989:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202998:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 202999:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203006:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203007:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203014:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203015:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203023:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203024:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203033:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203034:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203041:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203042:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203050:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203051:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203059:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203060:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203069:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203070:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203077:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203078:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203085:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203086:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203094:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203095:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203165:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203166:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203173:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203174:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203181:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203182:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203189:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203190:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203197:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203198:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203246:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203247:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203254:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203255:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203262:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203263:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203270:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203271:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203278:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203279:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203286:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203287:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203431:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203432:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203491:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203492:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203502:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203503:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203510:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203511:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203524:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203525:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203532:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203533:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203551:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203552:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203563:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203564:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203591:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203592:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203813:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203814:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203834:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 203835:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203898:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 203899:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {3{`RANDOM}};
  inflight = _RAND_13[95:0];
  _RAND_14 = {12{`RANDOM}};
  inflight_opcodes = _RAND_14[383:0];
  _RAND_15 = {12{`RANDOM}};
  inflight_sizes = _RAND_15[383:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {3{`RANDOM}};
  inflight_1 = _RAND_19[95:0];
  _RAND_20 = {12{`RANDOM}};
  inflight_sizes_1 = _RAND_20[383:0];
  _RAND_21 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  watchdog_1 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_22_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 203913:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 203914:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 203915:4]
  output        io_enq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  input         io_enq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  input  [2:0]  io_enq_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  input  [1:0]  io_enq_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  input  [6:0]  io_enq_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  input  [28:0] io_enq_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  input  [3:0]  io_enq_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  input  [31:0] io_enq_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  input         io_deq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  output        io_deq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  output [1:0]  io_deq_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  output [6:0]  io_deq_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  output [28:0] io_deq_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  output [3:0]  io_deq_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  output [31:0] io_deq_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 203916:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  reg [1:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  reg [6:0] ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [6:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [6:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  reg [28:0] ram_address [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [28:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [28:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  reg [3:0] ram_mask [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [3:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [3:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  reg [31:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [31:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire [31:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 203919:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 203920:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 203921:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.TinyRocketConfig.fir 203922:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.TinyRocketConfig.fir 203923:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.TinyRocketConfig.fir 203924:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.TinyRocketConfig.fir 203925:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 203926:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 203929:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 203944:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 203950:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.TinyRocketConfig.fir 203953:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.TinyRocketConfig.fir 203959:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.TinyRocketConfig.fir 203957:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 203969:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 203968:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 203967:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 203966:4]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 203965:4]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 203964:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 203963:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 203962:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 203918:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 203919:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 203919:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.TinyRocketConfig.fir 203932:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 203945:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 203920:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 203920:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.TinyRocketConfig.fir 203947:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 203951:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 203921:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 203921:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.TinyRocketConfig.fir 203954:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.TinyRocketConfig.fir 203955:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[28:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_16_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 204041:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 204042:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 204043:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [1:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [6:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [3:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [31:0] auto_in_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [1:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [6:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [31:0] auto_in_d_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [1:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [6:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [3:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output [31:0] auto_out_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [1:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [6:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
  input  [31:0] auto_out_d_bits_data // @[chipyard.TestHarness.TinyRocketConfig.fir 204044:4]
);
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire [1:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire [6:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire [1:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire [6:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [1:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [6:0] bundleOut_0_a_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [28:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [31:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire  bundleOut_0_a_q_io_enq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [1:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [6:0] bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [28:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire [31:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire  bundleOut_0_a_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire [1:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire [6:0] bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire [31:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire [6:0] bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire  bundleIn_0_d_q_io_deq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire [31:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
  TLMonitor_43_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 204051:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_22_inTestHarness bundleOut_0_a_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204078:4]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
  );
  Queue_5_inTestHarness bundleIn_0_d_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 204092:4]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Decoupled.scala 299:17 chipyard.TestHarness.TinyRocketConfig.fir 204090:4]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 204091:4]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 204091:4]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 204091:4]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 204091:4]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 204091:4]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 204091:4]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 204091:4]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 204091:4]
  assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 204091:4]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 Decoupled.scala 299:17 chipyard.TestHarness.TinyRocketConfig.fir 204104:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 204052:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 204053:4]
  assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Decoupled.scala 299:17 chipyard.TestHarness.TinyRocketConfig.fir 204090:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 204105:4]
  assign bundleOut_0_a_q_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 204079:4]
  assign bundleOut_0_a_q_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 204080:4]
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 204076:4]
  assign bundleIn_0_d_q_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 204093:4]
  assign bundleIn_0_d_q_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 204094:4]
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 204076:4]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 204076:4]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 204076:4]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 204076:4]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 204074:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 204076:4]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 204049:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 204077:4]
endmodule
module TLMonitor_44_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 204141:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 204142:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 204143:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input  [2:0]  io_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input  [1:0]  io_in_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input  [3:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input  [2:0]  io_in_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input  [1:0]  io_in_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input         io_in_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 204144:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 205589:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 205896:4]
  wire  _source_ok_T = io_in_a_bits_source == 2'h2; // @[Parameters.scala 46:9 chipyard.TestHarness.TinyRocketConfig.fir 204155:6]
  wire  _source_ok_T_1 = io_in_a_bits_source == 2'h1; // @[Parameters.scala 46:9 chipyard.TestHarness.TinyRocketConfig.fir 204156:6]
  wire  _source_ok_T_2 = io_in_a_bits_source == 2'h0; // @[Parameters.scala 46:9 chipyard.TestHarness.TinyRocketConfig.fir 204157:6]
  wire  _source_ok_T_3 = _source_ok_T | _source_ok_T_1; // @[Parameters.scala 1125:46 chipyard.TestHarness.TinyRocketConfig.fir 204163:6]
  wire  source_ok = _source_ok_T_3 | _source_ok_T_2; // @[Parameters.scala 1125:46 chipyard.TestHarness.TinyRocketConfig.fir 204164:6]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 204166:6]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 204168:6]
  wire [28:0] _GEN_71 = {{23'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.TinyRocketConfig.fir 204169:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.TinyRocketConfig.fir 204169:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.TinyRocketConfig.fir 204170:6]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49 chipyard.TestHarness.TinyRocketConfig.fir 204172:6]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.TinyRocketConfig.fir 204173:6]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81 chipyard.TestHarness.TinyRocketConfig.fir 204175:6]
  wire  _mask_T = io_in_a_bits_size >= 3'h2; // @[Misc.scala 205:21 chipyard.TestHarness.TinyRocketConfig.fir 204176:6]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 204177:6]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 204178:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 204179:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 204181:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 204182:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 204184:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 204185:6]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 204186:6]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 204187:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 204188:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 204189:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 204190:6]
  wire  mask_lo_lo = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 204191:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 204192:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 204193:6]
  wire  mask_lo_hi = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 204194:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 204195:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 204196:6]
  wire  mask_hi_lo = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 204197:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 204198:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 204199:6]
  wire  mask_hi_hi = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 204200:6]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 204203:6]
  wire  _T_33 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.TinyRocketConfig.fir 204237:6]
  wire [28:0] _T_45 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 204250:8]
  wire [29:0] _T_46 = {1'b0,$signed(_T_45)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 204251:8]
  wire [29:0] _T_48 = $signed(_T_46) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 204253:8]
  wire  _T_49 = $signed(_T_48) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 204254:8]
  wire  _T_55 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204260:8]
  wire  _T_72 = source_ok | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204285:8]
  wire  _T_73 = ~_T_72; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204286:8]
  wire  _T_76 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204293:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204294:8]
  wire  _T_79 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204300:8]
  wire  _T_80 = ~_T_79; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204301:8]
  wire  _T_81 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.TinyRocketConfig.fir 204306:8]
  wire  _T_83 = _T_81 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204308:8]
  wire  _T_84 = ~_T_83; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204309:8]
  wire [3:0] _T_85 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.TinyRocketConfig.fir 204314:8]
  wire  _T_86 = _T_85 == 4'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.TinyRocketConfig.fir 204315:8]
  wire  _T_88 = _T_86 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204317:8]
  wire  _T_89 = ~_T_88; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204318:8]
  wire  _T_90 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.TinyRocketConfig.fir 204323:8]
  wire  _T_92 = _T_90 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204325:8]
  wire  _T_93 = ~_T_92; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204326:8]
  wire  _T_94 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.TinyRocketConfig.fir 204332:6]
  wire  _T_146 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.TinyRocketConfig.fir 204409:8]
  wire  _T_148 = _T_146 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204411:8]
  wire  _T_149 = ~_T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204412:8]
  wire  _T_159 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.TinyRocketConfig.fir 204435:6]
  wire  _T_174 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.TinyRocketConfig.fir 204455:8]
  wire  _T_182 = _T_174 & _T_49; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 204463:8]
  wire  _T_185 = _T_182 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204466:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204467:8]
  wire  _T_193 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.TinyRocketConfig.fir 204486:8]
  wire  _T_195 = _T_193 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204488:8]
  wire  _T_196 = ~_T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204489:8]
  wire  _T_197 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.TinyRocketConfig.fir 204494:8]
  wire  _T_199 = _T_197 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204496:8]
  wire  _T_200 = ~_T_199; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204497:8]
  wire  _T_205 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.TinyRocketConfig.fir 204511:6]
  wire  _T_227 = source_ok & _T_182; // @[Monitor.scala 115:71 chipyard.TestHarness.TinyRocketConfig.fir 204534:8]
  wire  _T_229 = _T_227 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204536:8]
  wire  _T_230 = ~_T_229; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204537:8]
  wire  _T_245 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.TinyRocketConfig.fir 204573:6]
  wire [3:0] _T_281 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.TinyRocketConfig.fir 204626:8]
  wire [3:0] _T_282 = io_in_a_bits_mask & _T_281; // @[Monitor.scala 127:31 chipyard.TestHarness.TinyRocketConfig.fir 204627:8]
  wire  _T_283 = _T_282 == 4'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.TinyRocketConfig.fir 204628:8]
  wire  _T_285 = _T_283 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204630:8]
  wire  _T_286 = ~_T_285; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204631:8]
  wire  _T_287 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.TinyRocketConfig.fir 204637:6]
  wire  _T_316 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.TinyRocketConfig.fir 204679:8]
  wire  _T_318 = _T_316 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204681:8]
  wire  _T_319 = ~_T_318; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204682:8]
  wire  _T_324 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.TinyRocketConfig.fir 204696:6]
  wire  _T_353 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.TinyRocketConfig.fir 204738:8]
  wire  _T_355 = _T_353 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204740:8]
  wire  _T_356 = ~_T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204741:8]
  wire  _T_361 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.TinyRocketConfig.fir 204755:6]
  wire  _T_390 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.TinyRocketConfig.fir 204797:8]
  wire  _T_392 = _T_390 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204799:8]
  wire  _T_393 = ~_T_392; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204800:8]
  wire  _T_402 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.TinyRocketConfig.fir 204824:6]
  wire  _T_404 = _T_402 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204826:6]
  wire  _T_405 = ~_T_404; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204827:6]
  wire  _source_ok_T_4 = io_in_d_bits_source == 2'h2; // @[Parameters.scala 46:9 chipyard.TestHarness.TinyRocketConfig.fir 204832:6]
  wire  _source_ok_T_5 = io_in_d_bits_source == 2'h1; // @[Parameters.scala 46:9 chipyard.TestHarness.TinyRocketConfig.fir 204833:6]
  wire  _source_ok_T_6 = io_in_d_bits_source == 2'h0; // @[Parameters.scala 46:9 chipyard.TestHarness.TinyRocketConfig.fir 204834:6]
  wire  _source_ok_T_7 = _source_ok_T_4 | _source_ok_T_5; // @[Parameters.scala 1125:46 chipyard.TestHarness.TinyRocketConfig.fir 204840:6]
  wire  source_ok_1 = _source_ok_T_7 | _source_ok_T_6; // @[Parameters.scala 1125:46 chipyard.TestHarness.TinyRocketConfig.fir 204841:6]
  wire  _T_406 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.TinyRocketConfig.fir 204843:6]
  wire  _T_408 = source_ok_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204846:8]
  wire  _T_409 = ~_T_408; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204847:8]
  wire  _T_410 = io_in_d_bits_size >= 3'h2; // @[Monitor.scala 312:27 chipyard.TestHarness.TinyRocketConfig.fir 204852:8]
  wire  _T_412 = _T_410 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204854:8]
  wire  _T_413 = ~_T_412; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204855:8]
  wire  _T_414 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.TinyRocketConfig.fir 204860:8]
  wire  _T_416 = _T_414 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204862:8]
  wire  _T_417 = ~_T_416; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204863:8]
  wire  _T_418 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.TinyRocketConfig.fir 204868:8]
  wire  _T_420 = _T_418 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204870:8]
  wire  _T_421 = ~_T_420; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204871:8]
  wire  _T_422 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.TinyRocketConfig.fir 204876:8]
  wire  _T_424 = _T_422 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204878:8]
  wire  _T_425 = ~_T_424; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204879:8]
  wire  _T_426 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.TinyRocketConfig.fir 204885:6]
  wire  _T_437 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.TinyRocketConfig.fir 204909:8]
  wire  _T_439 = _T_437 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204911:8]
  wire  _T_440 = ~_T_439; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204912:8]
  wire  _T_441 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.TinyRocketConfig.fir 204917:8]
  wire  _T_443 = _T_441 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204919:8]
  wire  _T_444 = ~_T_443; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204920:8]
  wire  _T_454 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.TinyRocketConfig.fir 204943:6]
  wire  _T_474 = _T_422 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.TinyRocketConfig.fir 204984:8]
  wire  _T_476 = _T_474 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204986:8]
  wire  _T_477 = ~_T_476; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204987:8]
  wire  _T_483 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.TinyRocketConfig.fir 205002:6]
  wire  _T_500 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.TinyRocketConfig.fir 205037:6]
  wire  _T_518 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.TinyRocketConfig.fir 205073:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 205139:4]
  wire [3:0] a_first_beats1_decode = is_aligned_mask[5:2]; // @[Edges.scala 219:59 chipyard.TestHarness.TinyRocketConfig.fir 205144:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.TinyRocketConfig.fir 205146:4]
  reg [3:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205148:4]
  wire [3:0] a_first_counter1 = a_first_counter - 4'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 205150:4]
  wire  a_first = a_first_counter == 4'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 205151:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.TinyRocketConfig.fir 205162:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.TinyRocketConfig.fir 205163:4]
  reg [2:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.TinyRocketConfig.fir 205164:4]
  reg [1:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.TinyRocketConfig.fir 205165:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.TinyRocketConfig.fir 205166:4]
  wire  _T_547 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.TinyRocketConfig.fir 205167:4]
  wire  _T_548 = io_in_a_valid & _T_547; // @[Monitor.scala 389:19 chipyard.TestHarness.TinyRocketConfig.fir 205168:4]
  wire  _T_549 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.TinyRocketConfig.fir 205170:6]
  wire  _T_551 = _T_549 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205172:6]
  wire  _T_552 = ~_T_551; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205173:6]
  wire  _T_553 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.TinyRocketConfig.fir 205178:6]
  wire  _T_555 = _T_553 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205180:6]
  wire  _T_556 = ~_T_555; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205181:6]
  wire  _T_557 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.TinyRocketConfig.fir 205186:6]
  wire  _T_559 = _T_557 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205188:6]
  wire  _T_560 = ~_T_559; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205189:6]
  wire  _T_561 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.TinyRocketConfig.fir 205194:6]
  wire  _T_563 = _T_561 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205196:6]
  wire  _T_564 = ~_T_563; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205197:6]
  wire  _T_565 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.TinyRocketConfig.fir 205202:6]
  wire  _T_567 = _T_565 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205204:6]
  wire  _T_568 = ~_T_567; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205205:6]
  wire  _T_570 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.TinyRocketConfig.fir 205212:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 205220:4]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 205222:4]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 205224:4]
  wire [3:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:2]; // @[Edges.scala 219:59 chipyard.TestHarness.TinyRocketConfig.fir 205225:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.TinyRocketConfig.fir 205226:4]
  reg [3:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205228:4]
  wire [3:0] d_first_counter1 = d_first_counter - 4'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 205230:4]
  wire  d_first = d_first_counter == 4'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 205231:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.TinyRocketConfig.fir 205242:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.TinyRocketConfig.fir 205243:4]
  reg [2:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.TinyRocketConfig.fir 205244:4]
  reg [1:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.TinyRocketConfig.fir 205245:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.TinyRocketConfig.fir 205246:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.TinyRocketConfig.fir 205247:4]
  wire  _T_571 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.TinyRocketConfig.fir 205248:4]
  wire  _T_572 = io_in_d_valid & _T_571; // @[Monitor.scala 541:19 chipyard.TestHarness.TinyRocketConfig.fir 205249:4]
  wire  _T_573 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.TinyRocketConfig.fir 205251:6]
  wire  _T_575 = _T_573 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205253:6]
  wire  _T_576 = ~_T_575; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205254:6]
  wire  _T_577 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.TinyRocketConfig.fir 205259:6]
  wire  _T_579 = _T_577 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205261:6]
  wire  _T_580 = ~_T_579; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205262:6]
  wire  _T_581 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.TinyRocketConfig.fir 205267:6]
  wire  _T_583 = _T_581 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205269:6]
  wire  _T_584 = ~_T_583; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205270:6]
  wire  _T_585 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.TinyRocketConfig.fir 205275:6]
  wire  _T_587 = _T_585 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205277:6]
  wire  _T_588 = ~_T_587; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205278:6]
  wire  _T_589 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.TinyRocketConfig.fir 205283:6]
  wire  _T_591 = _T_589 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205285:6]
  wire  _T_592 = ~_T_591; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205286:6]
  wire  _T_593 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.TinyRocketConfig.fir 205291:6]
  wire  _T_595 = _T_593 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205293:6]
  wire  _T_596 = ~_T_595; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205294:6]
  wire  _T_598 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.TinyRocketConfig.fir 205301:4]
  reg [2:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 205310:4]
  reg [11:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 205311:4]
  reg [11:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 205312:4]
  reg [3:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205322:4]
  wire [3:0] a_first_counter1_1 = a_first_counter_1 - 4'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 205324:4]
  wire  a_first_1 = a_first_counter_1 == 4'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 205325:4]
  reg [3:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205344:4]
  wire [3:0] d_first_counter1_1 = d_first_counter_1 - 4'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 205346:4]
  wire  d_first_1 = d_first_counter_1 == 4'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 205347:4]
  wire [3:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.TinyRocketConfig.fir 205368:4]
  wire [4:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.TinyRocketConfig.fir 205368:4]
  wire [11:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.TinyRocketConfig.fir 205369:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.TinyRocketConfig.fir 205373:4]
  wire [15:0] _GEN_73 = {{4'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.TinyRocketConfig.fir 205374:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.TinyRocketConfig.fir 205374:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.TinyRocketConfig.fir 205375:4]
  wire [11:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.TinyRocketConfig.fir 205380:4]
  wire [15:0] _GEN_76 = {{4'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.TinyRocketConfig.fir 205385:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_76 & _a_opcode_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.TinyRocketConfig.fir 205385:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.TinyRocketConfig.fir 205386:4]
  wire  _T_599 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.TinyRocketConfig.fir 205410:4]
  wire [3:0] _a_set_wo_ready_T = 4'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.TinyRocketConfig.fir 205413:6]
  wire [3:0] _GEN_15 = _T_599 ? _a_set_wo_ready_T : 4'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.TinyRocketConfig.fir 205412:4 Monitor.scala 649:22 chipyard.TestHarness.TinyRocketConfig.fir 205414:6 chipyard.TestHarness.TinyRocketConfig.fir 205361:4]
  wire  _T_602 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.TinyRocketConfig.fir 205417:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.TinyRocketConfig.fir 205422:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.TinyRocketConfig.fir 205423:6]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.TinyRocketConfig.fir 205425:6]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.TinyRocketConfig.fir 205426:6]
  wire [3:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.TinyRocketConfig.fir 205428:6]
  wire [4:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.TinyRocketConfig.fir 205428:6]
  wire [3:0] a_opcodes_set_interm = _T_602 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 205419:4 Monitor.scala 654:28 chipyard.TestHarness.TinyRocketConfig.fir 205424:6 chipyard.TestHarness.TinyRocketConfig.fir 205407:4]
  wire [34:0] _GEN_79 = {{31'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.TinyRocketConfig.fir 205429:6]
  wire [34:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.TinyRocketConfig.fir 205429:6]
  wire [3:0] a_sizes_set_interm = _T_602 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 205419:4 Monitor.scala 655:28 chipyard.TestHarness.TinyRocketConfig.fir 205427:6 chipyard.TestHarness.TinyRocketConfig.fir 205409:4]
  wire [34:0] _GEN_81 = {{31'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.TinyRocketConfig.fir 205432:6]
  wire [34:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.TinyRocketConfig.fir 205432:6]
  wire [2:0] _T_604 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.TinyRocketConfig.fir 205434:6]
  wire  _T_606 = ~_T_604[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.TinyRocketConfig.fir 205436:6]
  wire  _T_608 = _T_606 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205438:6]
  wire  _T_609 = ~_T_608; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205439:6]
  wire [3:0] _GEN_16 = _T_602 ? _a_set_wo_ready_T : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 205419:4 Monitor.scala 653:28 chipyard.TestHarness.TinyRocketConfig.fir 205421:6 chipyard.TestHarness.TinyRocketConfig.fir 205359:4]
  wire [34:0] _GEN_19 = _T_602 ? _a_opcodes_set_T_1 : 35'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 205419:4 Monitor.scala 656:28 chipyard.TestHarness.TinyRocketConfig.fir 205430:6 chipyard.TestHarness.TinyRocketConfig.fir 205363:4]
  wire [34:0] _GEN_20 = _T_602 ? _a_sizes_set_T_1 : 35'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 205419:4 Monitor.scala 657:28 chipyard.TestHarness.TinyRocketConfig.fir 205433:6 chipyard.TestHarness.TinyRocketConfig.fir 205365:4]
  wire  _T_610 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.TinyRocketConfig.fir 205454:4]
  wire  _T_612 = ~_T_406; // @[Monitor.scala 671:74 chipyard.TestHarness.TinyRocketConfig.fir 205456:4]
  wire  _T_613 = _T_610 & _T_612; // @[Monitor.scala 671:71 chipyard.TestHarness.TinyRocketConfig.fir 205457:4]
  wire [3:0] _d_clr_wo_ready_T = 4'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.TinyRocketConfig.fir 205459:6]
  wire [3:0] _GEN_21 = _T_613 ? _d_clr_wo_ready_T : 4'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.TinyRocketConfig.fir 205458:4 Monitor.scala 672:22 chipyard.TestHarness.TinyRocketConfig.fir 205460:6 chipyard.TestHarness.TinyRocketConfig.fir 205448:4]
  wire  _T_615 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.TinyRocketConfig.fir 205463:4]
  wire  _T_618 = _T_615 & _T_612; // @[Monitor.scala 675:72 chipyard.TestHarness.TinyRocketConfig.fir 205466:4]
  wire [46:0] _GEN_83 = {{31'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.TinyRocketConfig.fir 205475:6]
  wire [46:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.TinyRocketConfig.fir 205475:6]
  wire [3:0] _GEN_22 = _T_618 ? _d_clr_wo_ready_T : 4'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 205467:4 Monitor.scala 676:21 chipyard.TestHarness.TinyRocketConfig.fir 205469:6 chipyard.TestHarness.TinyRocketConfig.fir 205446:4]
  wire [46:0] _GEN_23 = _T_618 ? _d_opcodes_clr_T_5 : 47'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 205467:4 Monitor.scala 677:21 chipyard.TestHarness.TinyRocketConfig.fir 205476:6 chipyard.TestHarness.TinyRocketConfig.fir 205450:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.TinyRocketConfig.fir 205492:6]
  wire  same_cycle_resp = _T_599 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.TinyRocketConfig.fir 205493:6]
  wire [2:0] _T_623 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.TinyRocketConfig.fir 205494:6]
  wire  _T_625 = _T_623[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.TinyRocketConfig.fir 205496:6]
  wire  _T_627 = _T_625 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205498:6]
  wire  _T_628 = ~_T_627; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205499:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8]
  wire  _T_629 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 205505:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 205506:8 Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 205506:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 205506:8 Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 205506:8]
  wire  _T_630 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 205506:8]
  wire  _T_631 = _T_629 | _T_630; // @[Monitor.scala 685:77 chipyard.TestHarness.TinyRocketConfig.fir 205507:8]
  wire  _T_633 = _T_631 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205509:8]
  wire  _T_634 = ~_T_633; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205510:8]
  wire  _T_635 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.TinyRocketConfig.fir 205515:8]
  wire  _T_637 = _T_635 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205517:8]
  wire  _T_638 = ~_T_637; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205518:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205366:4 Monitor.scala 634:21 chipyard.TestHarness.TinyRocketConfig.fir 205376:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8]
  wire  _T_640 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 205526:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 205528:8 Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 205528:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 205528:8 Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 205528:8]
  wire  _T_642 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 205528:8]
  wire  _T_643 = _T_640 | _T_642; // @[Monitor.scala 689:72 chipyard.TestHarness.TinyRocketConfig.fir 205529:8]
  wire  _T_645 = _T_643 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205531:8]
  wire  _T_646 = ~_T_645; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205532:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205377:4 Monitor.scala 638:19 chipyard.TestHarness.TinyRocketConfig.fir 205387:4]
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.TinyRocketConfig.fir 205537:8]
  wire  _T_647 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.TinyRocketConfig.fir 205537:8]
  wire  _T_649 = _T_647 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205539:8]
  wire  _T_650 = ~_T_649; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205540:8]
  wire  _T_652 = _T_610 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.TinyRocketConfig.fir 205548:4]
  wire  _T_653 = _T_652 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.TinyRocketConfig.fir 205549:4]
  wire  _T_655 = _T_653 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.TinyRocketConfig.fir 205551:4]
  wire  _T_657 = _T_655 & _T_612; // @[Monitor.scala 694:116 chipyard.TestHarness.TinyRocketConfig.fir 205553:4]
  wire  _T_658 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.TinyRocketConfig.fir 205555:6]
  wire  _T_659 = _T_658 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.TinyRocketConfig.fir 205556:6]
  wire  _T_661 = _T_659 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205558:6]
  wire  _T_662 = ~_T_661; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205559:6]
  wire [2:0] a_set_wo_ready = _GEN_15[2:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205360:4]
  wire [2:0] d_clr_wo_ready = _GEN_21[2:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205447:4]
  wire  _T_663 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.TinyRocketConfig.fir 205565:4]
  wire  _T_664 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.TinyRocketConfig.fir 205566:4]
  wire  _T_665 = ~_T_664; // @[Monitor.scala 699:51 chipyard.TestHarness.TinyRocketConfig.fir 205567:4]
  wire  _T_666 = _T_663 | _T_665; // @[Monitor.scala 699:48 chipyard.TestHarness.TinyRocketConfig.fir 205568:4]
  wire  _T_668 = _T_666 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205570:4]
  wire  _T_669 = ~_T_668; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205571:4]
  wire [2:0] a_set = _GEN_16[2:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205358:4]
  wire [2:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.TinyRocketConfig.fir 205576:4]
  wire [2:0] d_clr = _GEN_22[2:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205445:4]
  wire [2:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.TinyRocketConfig.fir 205577:4]
  wire [2:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.TinyRocketConfig.fir 205578:4]
  wire [11:0] a_opcodes_set = _GEN_19[11:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205362:4]
  wire [11:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.TinyRocketConfig.fir 205580:4]
  wire [11:0] d_opcodes_clr = _GEN_23[11:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205449:4]
  wire [11:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.TinyRocketConfig.fir 205581:4]
  wire [11:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.TinyRocketConfig.fir 205582:4]
  wire [11:0] a_sizes_set = _GEN_20[11:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205364:4]
  wire [11:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.TinyRocketConfig.fir 205584:4]
  wire [11:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.TinyRocketConfig.fir 205586:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 205588:4]
  wire  _T_670 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.TinyRocketConfig.fir 205591:4]
  wire  _T_671 = ~_T_670; // @[Monitor.scala 709:16 chipyard.TestHarness.TinyRocketConfig.fir 205592:4]
  wire  _T_672 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.TinyRocketConfig.fir 205593:4]
  wire  _T_673 = _T_671 | _T_672; // @[Monitor.scala 709:30 chipyard.TestHarness.TinyRocketConfig.fir 205594:4]
  wire  _T_674 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.TinyRocketConfig.fir 205595:4]
  wire  _T_675 = _T_673 | _T_674; // @[Monitor.scala 709:47 chipyard.TestHarness.TinyRocketConfig.fir 205596:4]
  wire  _T_677 = _T_675 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205598:4]
  wire  _T_678 = ~_T_677; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205599:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.TinyRocketConfig.fir 205605:4]
  wire  _T_681 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.TinyRocketConfig.fir 205609:4]
  reg [2:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.TinyRocketConfig.fir 205613:4]
  reg [11:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 205615:4]
  reg [3:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205650:4]
  wire [3:0] d_first_counter1_2 = d_first_counter_2 - 4'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 205652:4]
  wire  d_first_2 = d_first_counter_2 == 4'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 205653:4]
  wire [11:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.TinyRocketConfig.fir 205686:4]
  wire [15:0] _GEN_91 = {{4'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.TinyRocketConfig.fir 205691:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_91 & _a_opcode_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.TinyRocketConfig.fir 205691:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.TinyRocketConfig.fir 205692:4]
  wire  _T_699 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.TinyRocketConfig.fir 205770:4]
  wire  _T_701 = _T_699 & _T_406; // @[Monitor.scala 779:71 chipyard.TestHarness.TinyRocketConfig.fir 205772:4]
  wire  _T_703 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.TinyRocketConfig.fir 205778:4]
  wire  _T_705 = _T_703 & _T_406; // @[Monitor.scala 783:72 chipyard.TestHarness.TinyRocketConfig.fir 205780:4]
  wire [3:0] _GEN_67 = _T_705 ? _d_clr_wo_ready_T : 4'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.TinyRocketConfig.fir 205781:4 Monitor.scala 784:21 chipyard.TestHarness.TinyRocketConfig.fir 205783:6 chipyard.TestHarness.TinyRocketConfig.fir 205762:4]
  wire [46:0] _GEN_68 = _T_705 ? _d_opcodes_clr_T_5 : 47'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.TinyRocketConfig.fir 205781:4 Monitor.scala 785:21 chipyard.TestHarness.TinyRocketConfig.fir 205790:6 chipyard.TestHarness.TinyRocketConfig.fir 205766:4]
  wire [2:0] _T_709 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.TinyRocketConfig.fir 205816:6]
  wire  _T_713 = _T_709[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205820:6]
  wire  _T_714 = ~_T_713; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205821:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205674:4 Monitor.scala 747:21 chipyard.TestHarness.TinyRocketConfig.fir 205693:4]
  wire  _T_719 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.TinyRocketConfig.fir 205839:8]
  wire  _T_721 = _T_719 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205841:8]
  wire  _T_722 = ~_T_721; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205842:8]
  wire [2:0] d_clr_1 = _GEN_67[2:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205761:4]
  wire [2:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.TinyRocketConfig.fir 205884:4]
  wire [2:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.TinyRocketConfig.fir 205885:4]
  wire [11:0] d_opcodes_clr_1 = _GEN_68[11:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 205765:4]
  wire [11:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.TinyRocketConfig.fir 205888:4]
  wire [11:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.TinyRocketConfig.fir 205893:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.TinyRocketConfig.fir 205895:4]
  wire  _T_739 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.TinyRocketConfig.fir 205898:4]
  wire  _T_740 = ~_T_739; // @[Monitor.scala 816:16 chipyard.TestHarness.TinyRocketConfig.fir 205899:4]
  wire  _T_741 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.TinyRocketConfig.fir 205900:4]
  wire  _T_742 = _T_740 | _T_741; // @[Monitor.scala 816:30 chipyard.TestHarness.TinyRocketConfig.fir 205901:4]
  wire  _T_743 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.TinyRocketConfig.fir 205902:4]
  wire  _T_744 = _T_742 | _T_743; // @[Monitor.scala 816:47 chipyard.TestHarness.TinyRocketConfig.fir 205903:4]
  wire  _T_746 = _T_744 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205905:4]
  wire  _T_747 = ~_T_746; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205906:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.TinyRocketConfig.fir 205912:4]
  wire  _GEN_98 = io_in_a_valid & _T_33; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204262:10]
  wire  _GEN_114 = io_in_a_valid & _T_94; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204357:10]
  wire  _GEN_132 = io_in_a_valid & _T_159; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204451:10]
  wire  _GEN_146 = io_in_a_valid & _T_205; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204539:10]
  wire  _GEN_156 = io_in_a_valid & _T_245; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204601:10]
  wire  _GEN_166 = io_in_a_valid & _T_287; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204662:10]
  wire  _GEN_176 = io_in_a_valid & _T_324; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204721:10]
  wire  _GEN_186 = io_in_a_valid & _T_361; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204780:10]
  wire  _GEN_198 = io_in_d_valid & _T_406; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204849:10]
  wire  _GEN_208 = io_in_d_valid & _T_426; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204891:10]
  wire  _GEN_222 = io_in_d_valid & _T_454; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204949:10]
  wire  _GEN_236 = io_in_d_valid & _T_483; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205008:10]
  wire  _GEN_244 = io_in_d_valid & _T_500; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205043:10]
  wire  _GEN_252 = io_in_d_valid & _T_518; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205079:10]
  wire  _GEN_260 = _T_613 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205512:10]
  wire  _GEN_265 = _T_613 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205534:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 205589:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 205896:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205148:4]
      a_first_counter <= 4'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205148:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 205158:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 205159:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 205147:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 4'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_570) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 205213:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.TinyRocketConfig.fir 205214:6]
    end
    if (_T_570) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 205213:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.TinyRocketConfig.fir 205215:6]
    end
    if (_T_570) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 205213:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.TinyRocketConfig.fir 205216:6]
    end
    if (_T_570) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 205213:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.TinyRocketConfig.fir 205217:6]
    end
    if (_T_570) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 205213:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.TinyRocketConfig.fir 205218:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205228:4]
      d_first_counter <= 4'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205228:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 205238:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 205239:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 205227:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 4'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_598) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 205302:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.TinyRocketConfig.fir 205303:6]
    end
    if (_T_598) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 205302:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.TinyRocketConfig.fir 205304:6]
    end
    if (_T_598) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 205302:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.TinyRocketConfig.fir 205305:6]
    end
    if (_T_598) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 205302:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.TinyRocketConfig.fir 205306:6]
    end
    if (_T_598) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 205302:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.TinyRocketConfig.fir 205307:6]
    end
    if (_T_598) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 205302:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.TinyRocketConfig.fir 205308:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 205310:4]
      inflight <= 3'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 205310:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.TinyRocketConfig.fir 205579:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 205311:4]
      inflight_opcodes <= 12'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 205311:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.TinyRocketConfig.fir 205583:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 205312:4]
      inflight_sizes <= 12'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 205312:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.TinyRocketConfig.fir 205587:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205322:4]
      a_first_counter_1 <= 4'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205322:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 205332:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 205333:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 205147:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 4'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205344:4]
      d_first_counter_1 <= 4'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205344:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 205354:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 205355:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 205227:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 4'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 205588:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 205588:4]
    end else if (_T_681) begin // @[Monitor.scala 712:47 chipyard.TestHarness.TinyRocketConfig.fir 205610:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.TinyRocketConfig.fir 205611:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.TinyRocketConfig.fir 205606:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.TinyRocketConfig.fir 205613:4]
      inflight_1 <= 3'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.TinyRocketConfig.fir 205613:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.TinyRocketConfig.fir 205886:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 205615:4]
      inflight_sizes_1 <= 12'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 205615:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.TinyRocketConfig.fir 205894:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205650:4]
      d_first_counter_2 <= 4'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 205650:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 205660:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 205661:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 205227:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 4'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.TinyRocketConfig.fir 205895:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.TinyRocketConfig.fir 205895:4]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47 chipyard.TestHarness.TinyRocketConfig.fir 205919:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.TinyRocketConfig.fir 205920:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.TinyRocketConfig.fir 205913:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_33 & _T_55) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204262:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_55) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204263:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_55) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204281:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_55) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204282:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_73) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204288:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_73) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204289:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204296:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204297:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_80) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204303:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_80) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204304:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204311:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204312:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_89) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204320:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_89) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204321:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_93) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204328:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_93) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204329:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_94 & _T_55) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204357:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_55) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204358:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_55) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204376:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_55) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204377:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_73) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204383:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_73) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204384:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204391:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204392:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_80) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204398:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_80) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204399:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204406:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204407:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_149) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204414:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_149) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204415:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_89) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204423:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_89) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204424:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_93) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204431:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_93) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204432:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_159 & _T_73) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204451:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_73) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204452:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204469:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204470:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_73) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204476:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_73) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204477:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_80) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204483:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_80) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204484:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_196) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204491:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_196) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204492:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_200) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204499:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_200) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204500:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_93) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204507:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_93) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204508:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_205 & _T_230) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204539:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_230) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204540:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_73) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204546:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_73) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204547:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_80) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204553:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_80) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204554:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_196) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204561:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_196) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204562:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_200) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204569:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_200) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204570:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_245 & _T_230) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204601:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_230) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204602:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_73) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204608:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_73) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204609:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_80) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204615:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_80) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204616:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_196) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204623:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_196) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204624:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_286) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204633:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_286) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204634:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_287 & _T_55) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204662:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_55) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204663:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_73) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204669:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_73) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204670:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_80) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204676:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_80) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204677:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_319) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204684:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_319) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204685:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_200) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204692:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_200) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204693:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_324 & _T_55) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204721:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_55) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204722:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_73) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204728:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_73) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204729:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_80) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204735:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_80) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204736:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_356) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204743:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_356) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204744:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_200) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204751:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_200) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204752:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_361 & _T_55) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204780:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_55) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204781:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_73) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204787:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_73) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204788:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_80) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204794:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_80) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204795:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_393) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204802:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_393) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204803:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_200) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204810:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_200) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204811:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_93) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204818:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_93) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 204819:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_405) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204829:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_405) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204830:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_406 & _T_409) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204849:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_409) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204850:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_413) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204857:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_413) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204858:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204865:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_417) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204866:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204873:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_421) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204874:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_425) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204881:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_425) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204882:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_426 & _T_409) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204891:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_409) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204892:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_55) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204898:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_55) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204899:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_413) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204906:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_413) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204907:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_440) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204914:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_440) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204915:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_444) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204922:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_444) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204923:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204930:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_421) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204931:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_425) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204939:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_425) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204940:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_454 & _T_409) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204949:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_409) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204950:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_55) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204956:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_55) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204957:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_413) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204964:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_413) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204965:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_440) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204972:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_440) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204973:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_444) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204980:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_444) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204981:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_477) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204989:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_477) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204990:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_425) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204998:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_425) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 204999:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_483 & _T_409) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205008:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_409) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205009:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205016:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_417) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205017:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205024:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_421) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205025:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_425) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205033:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_425) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205034:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_500 & _T_409) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205043:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_409) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205044:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205051:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_417) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205052:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_477) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205060:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_477) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205061:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_425) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205069:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_425) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205070:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_518 & _T_409) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205079:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_409) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205080:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205087:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_417) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205088:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205095:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_421) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205096:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_425) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205104:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_425) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205105:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_548 & _T_552) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205175:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_548 & _T_552) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205176:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_548 & _T_556) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205183:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_548 & _T_556) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205184:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_548 & _T_560) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205191:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_548 & _T_560) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205192:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_548 & _T_564) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205199:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_548 & _T_564) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205200:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_548 & _T_568) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205207:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_548 & _T_568) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205208:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_572 & _T_576) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205256:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_572 & _T_576) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205257:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_572 & _T_580) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205264:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_572 & _T_580) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205265:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_572 & _T_584) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205272:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_572 & _T_584) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205273:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_572 & _T_588) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205280:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_572 & _T_588) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205281:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_572 & _T_592) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205288:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_572 & _T_592) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205289:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_572 & _T_596) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205296:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_572 & _T_596) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205297:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_602 & _T_609) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205441:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_602 & _T_609) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205442:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_613 & _T_628) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205501:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_613 & _T_628) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205502:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_613 & same_cycle_resp & _T_634) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205512:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_634) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205513:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_638) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205520:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_638) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205521:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_613 & ~same_cycle_resp & _T_646) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205534:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_646) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205535:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & _T_650) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205542:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_650) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205543:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_657 & _T_662) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205561:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_657 & _T_662) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205562:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_669) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205573:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_669) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205574:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_678) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205601:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_678) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205602:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_701 & _T_714) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205823:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_701 & _T_714) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205824:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_701 & _T_722) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205844:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_701 & _T_722) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 205845:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_747) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205908:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_747) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 205909:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  inflight_opcodes = _RAND_14[11:0];
  _RAND_15 = {1{`RANDOM}};
  inflight_sizes = _RAND_15[11:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_1 = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_20[11:0];
  _RAND_21 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  watchdog_1 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater_7_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 205923:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 205924:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 205925:4]
  input         io_repeat, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  output        io_full, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  output        io_enq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  input         io_enq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  input  [2:0]  io_enq_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  input  [2:0]  io_enq_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  input  [1:0]  io_enq_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  input  [28:0] io_enq_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  input  [3:0]  io_enq_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  input         io_deq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  output        io_deq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  output [2:0]  io_deq_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  output [1:0]  io_deq_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  output [28:0] io_deq_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  output [3:0]  io_deq_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 205926:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21 chipyard.TestHarness.TinyRocketConfig.fir 205928:4]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18 chipyard.TestHarness.TinyRocketConfig.fir 205929:4]
  reg [2:0] saved_param; // @[Repeater.scala 20:18 chipyard.TestHarness.TinyRocketConfig.fir 205929:4]
  reg [2:0] saved_size; // @[Repeater.scala 20:18 chipyard.TestHarness.TinyRocketConfig.fir 205929:4]
  reg [1:0] saved_source; // @[Repeater.scala 20:18 chipyard.TestHarness.TinyRocketConfig.fir 205929:4]
  reg [28:0] saved_address; // @[Repeater.scala 20:18 chipyard.TestHarness.TinyRocketConfig.fir 205929:4]
  reg [3:0] saved_mask; // @[Repeater.scala 20:18 chipyard.TestHarness.TinyRocketConfig.fir 205929:4]
  reg  saved_corrupt; // @[Repeater.scala 20:18 chipyard.TestHarness.TinyRocketConfig.fir 205929:4]
  wire  _io_enq_ready_T = ~full; // @[Repeater.scala 24:35 chipyard.TestHarness.TinyRocketConfig.fir 205932:4]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 205945:4]
  wire  _T_1 = _T & io_repeat; // @[Repeater.scala 28:23 chipyard.TestHarness.TinyRocketConfig.fir 205946:4]
  wire  _GEN_0 = _T_1 | full; // @[Repeater.scala 28:38 chipyard.TestHarness.TinyRocketConfig.fir 205947:4 Repeater.scala 28:45 chipyard.TestHarness.TinyRocketConfig.fir 205948:6 Repeater.scala 19:21 chipyard.TestHarness.TinyRocketConfig.fir 205928:4]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 205958:4]
  wire  _T_3 = ~io_repeat; // @[Repeater.scala 29:26 chipyard.TestHarness.TinyRocketConfig.fir 205959:4]
  wire  _T_4 = _T_2 & _T_3; // @[Repeater.scala 29:23 chipyard.TestHarness.TinyRocketConfig.fir 205960:4]
  assign io_full = full; // @[Repeater.scala 26:11 chipyard.TestHarness.TinyRocketConfig.fir 205944:4]
  assign io_enq_ready = io_deq_ready & _io_enq_ready_T; // @[Repeater.scala 24:32 chipyard.TestHarness.TinyRocketConfig.fir 205933:4]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32 chipyard.TestHarness.TinyRocketConfig.fir 205930:4]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21 chipyard.TestHarness.TinyRocketConfig.fir 205935:4]
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; // @[Repeater.scala 25:21 chipyard.TestHarness.TinyRocketConfig.fir 205935:4]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21 chipyard.TestHarness.TinyRocketConfig.fir 205935:4]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21 chipyard.TestHarness.TinyRocketConfig.fir 205935:4]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21 chipyard.TestHarness.TinyRocketConfig.fir 205935:4]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21 chipyard.TestHarness.TinyRocketConfig.fir 205935:4]
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; // @[Repeater.scala 25:21 chipyard.TestHarness.TinyRocketConfig.fir 205935:4]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21 chipyard.TestHarness.TinyRocketConfig.fir 205928:4]
      full <= 1'h0; // @[Repeater.scala 19:21 chipyard.TestHarness.TinyRocketConfig.fir 205928:4]
    end else if (_T_4) begin // @[Repeater.scala 29:38 chipyard.TestHarness.TinyRocketConfig.fir 205961:4]
      full <= 1'h0; // @[Repeater.scala 29:45 chipyard.TestHarness.TinyRocketConfig.fir 205962:6]
    end else begin
      full <= _GEN_0;
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.TinyRocketConfig.fir 205947:4]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62 chipyard.TestHarness.TinyRocketConfig.fir 205956:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.TinyRocketConfig.fir 205947:4]
      saved_param <= io_enq_bits_param; // @[Repeater.scala 28:62 chipyard.TestHarness.TinyRocketConfig.fir 205955:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.TinyRocketConfig.fir 205947:4]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62 chipyard.TestHarness.TinyRocketConfig.fir 205954:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.TinyRocketConfig.fir 205947:4]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62 chipyard.TestHarness.TinyRocketConfig.fir 205953:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.TinyRocketConfig.fir 205947:4]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62 chipyard.TestHarness.TinyRocketConfig.fir 205952:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.TinyRocketConfig.fir 205947:4]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62 chipyard.TestHarness.TinyRocketConfig.fir 205951:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.TinyRocketConfig.fir 205947:4]
      saved_corrupt <= io_enq_bits_corrupt; // @[Repeater.scala 28:62 chipyard.TestHarness.TinyRocketConfig.fir 205949:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  saved_address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  saved_mask = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  saved_corrupt = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter_8_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 205965:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 205966:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 205967:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [2:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [1:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [3:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [31:0] auto_in_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [2:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [1:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [31:0] auto_in_d_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [1:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [6:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [3:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output [31:0] auto_out_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [1:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [6:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input         auto_out_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input  [31:0] auto_out_d_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 205968:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire [1:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire [1:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
  wire  repeater_clock; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire  repeater_reset; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [2:0] repeater_io_enq_bits_opcode; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [2:0] repeater_io_enq_bits_param; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [1:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [28:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [3:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire  repeater_io_enq_bits_corrupt; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [2:0] repeater_io_deq_bits_opcode; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [2:0] repeater_io_deq_bits_param; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [1:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [28:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire [3:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  wire  repeater_io_deq_bits_corrupt; // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
  reg [3:0] acknum; // @[Fragmenter.scala 189:29 chipyard.TestHarness.TinyRocketConfig.fir 206002:4]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24 chipyard.TestHarness.TinyRocketConfig.fir 206003:4]
  reg  dToggle; // @[Fragmenter.scala 191:30 chipyard.TestHarness.TinyRocketConfig.fir 206004:4]
  wire [3:0] dFragnum = auto_out_d_bits_source[3:0]; // @[Fragmenter.scala 192:41 chipyard.TestHarness.TinyRocketConfig.fir 206005:4]
  wire  dFirst = acknum == 4'h0; // @[Fragmenter.scala 193:29 chipyard.TestHarness.TinyRocketConfig.fir 206006:4]
  wire  dLast = dFragnum == 4'h0; // @[Fragmenter.scala 194:30 chipyard.TestHarness.TinyRocketConfig.fir 206007:4]
  wire [3:0] _dsizeOH_T = 4'h1 << auto_out_d_bits_size; // @[OneHot.scala 65:12 chipyard.TestHarness.TinyRocketConfig.fir 206009:4]
  wire [2:0] dsizeOH = _dsizeOH_T[2:0]; // @[OneHot.scala 65:27 chipyard.TestHarness.TinyRocketConfig.fir 206010:4]
  wire [4:0] _dsizeOH1_T_1 = 5'h3 << auto_out_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 206012:4]
  wire [1:0] dsizeOH1 = ~_dsizeOH1_T_1[1:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 206014:4]
  wire  dHasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.TinyRocketConfig.fir 206015:4]
  wire  ack_decrement = dHasData | dsizeOH[2]; // @[Fragmenter.scala 204:32 chipyard.TestHarness.TinyRocketConfig.fir 206032:4]
  wire [5:0] _dFirst_size_T = {dFragnum, 2'h0}; // @[Fragmenter.scala 206:47 chipyard.TestHarness.TinyRocketConfig.fir 206033:4]
  wire [5:0] _GEN_7 = {{4'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69 chipyard.TestHarness.TinyRocketConfig.fir 206034:4]
  wire [5:0] dFirst_size_lo = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69 chipyard.TestHarness.TinyRocketConfig.fir 206034:4]
  wire [6:0] _dFirst_size_T_1 = {dFirst_size_lo, 1'h0}; // @[package.scala 232:35 chipyard.TestHarness.TinyRocketConfig.fir 206035:4]
  wire [6:0] _dFirst_size_T_2 = _dFirst_size_T_1 | 7'h1; // @[package.scala 232:40 chipyard.TestHarness.TinyRocketConfig.fir 206036:4]
  wire [6:0] _dFirst_size_T_3 = {1'h0,dFirst_size_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 206037:4]
  wire [6:0] _dFirst_size_T_4 = ~_dFirst_size_T_3; // @[package.scala 232:53 chipyard.TestHarness.TinyRocketConfig.fir 206038:4]
  wire [6:0] _dFirst_size_T_5 = _dFirst_size_T_2 & _dFirst_size_T_4; // @[package.scala 232:51 chipyard.TestHarness.TinyRocketConfig.fir 206039:4]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_5[6:4]; // @[OneHot.scala 30:18 chipyard.TestHarness.TinyRocketConfig.fir 206040:4]
  wire [3:0] dFirst_size_lo_1 = _dFirst_size_T_5[3:0]; // @[OneHot.scala 31:18 chipyard.TestHarness.TinyRocketConfig.fir 206041:4]
  wire  dFirst_size_hi_1 = |dFirst_size_hi; // @[OneHot.scala 32:14 chipyard.TestHarness.TinyRocketConfig.fir 206042:4]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28 chipyard.TestHarness.TinyRocketConfig.fir 206043:4]
  wire [3:0] _dFirst_size_T_6 = _GEN_8 | dFirst_size_lo_1; // @[OneHot.scala 32:28 chipyard.TestHarness.TinyRocketConfig.fir 206043:4]
  wire [1:0] dFirst_size_hi_2 = _dFirst_size_T_6[3:2]; // @[OneHot.scala 30:18 chipyard.TestHarness.TinyRocketConfig.fir 206044:4]
  wire [1:0] dFirst_size_lo_2 = _dFirst_size_T_6[1:0]; // @[OneHot.scala 31:18 chipyard.TestHarness.TinyRocketConfig.fir 206045:4]
  wire  dFirst_size_hi_3 = |dFirst_size_hi_2; // @[OneHot.scala 32:14 chipyard.TestHarness.TinyRocketConfig.fir 206046:4]
  wire [1:0] _dFirst_size_T_7 = dFirst_size_hi_2 | dFirst_size_lo_2; // @[OneHot.scala 32:28 chipyard.TestHarness.TinyRocketConfig.fir 206047:4]
  wire  dFirst_size_lo_3 = _dFirst_size_T_7[1]; // @[CircuitMath.scala 30:8 chipyard.TestHarness.TinyRocketConfig.fir 206048:4]
  wire [2:0] dFirst_size = {dFirst_size_hi_1,dFirst_size_hi_3,dFirst_size_lo_3}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 206050:4]
  wire  _drop_T = ~dHasData; // @[Fragmenter.scala 222:20 chipyard.TestHarness.TinyRocketConfig.fir 206063:4]
  wire  _drop_T_2 = ~dLast; // @[Fragmenter.scala 222:33 chipyard.TestHarness.TinyRocketConfig.fir 206065:4]
  wire  drop = _drop_T & _drop_T_2; // @[Fragmenter.scala 222:30 chipyard.TestHarness.TinyRocketConfig.fir 206066:4]
  wire  bundleOut_0_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35 chipyard.TestHarness.TinyRocketConfig.fir 206067:4]
  wire  _T_7 = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 206051:4]
  wire [3:0] _GEN_9 = {{3'd0}, ack_decrement}; // @[Fragmenter.scala 209:55 chipyard.TestHarness.TinyRocketConfig.fir 206053:6]
  wire [3:0] _acknum_T_1 = acknum - _GEN_9; // @[Fragmenter.scala 209:55 chipyard.TestHarness.TinyRocketConfig.fir 206054:6]
  wire  _bundleIn_0_d_valid_T = ~drop; // @[Fragmenter.scala 224:39 chipyard.TestHarness.TinyRocketConfig.fir 206069:4]
  wire  _aFrag_T = repeater_io_deq_bits_size > 3'h2; // @[Fragmenter.scala 285:31 chipyard.TestHarness.TinyRocketConfig.fir 206102:4]
  wire [2:0] aFrag = _aFrag_T ? 3'h2 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24 chipyard.TestHarness.TinyRocketConfig.fir 206103:4]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 206105:4]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 206107:4]
  wire [8:0] _aFragOH1_T_1 = 9'h3 << aFrag; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 206109:4]
  wire [1:0] aFragOH1 = ~_aFragOH1_T_1[1:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 206111:4]
  wire  aHasData = ~repeater_io_deq_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.TinyRocketConfig.fir 206113:4]
  reg [3:0] gennum; // @[Fragmenter.scala 291:29 chipyard.TestHarness.TinyRocketConfig.fir 206115:4]
  wire  aFirst = gennum == 4'h0; // @[Fragmenter.scala 292:29 chipyard.TestHarness.TinyRocketConfig.fir 206116:4]
  wire [3:0] _old_gennum1_T_2 = gennum - 4'h1; // @[Fragmenter.scala 293:79 chipyard.TestHarness.TinyRocketConfig.fir 206119:4]
  wire [3:0] old_gennum1 = aFirst ? aOrigOH1[5:2] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30 chipyard.TestHarness.TinyRocketConfig.fir 206120:4]
  wire [3:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28 chipyard.TestHarness.TinyRocketConfig.fir 206121:4]
  wire [3:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26 chipyard.TestHarness.TinyRocketConfig.fir 206124:4]
  reg  aToggle_r; // @[Reg.scala 15:16 chipyard.TestHarness.TinyRocketConfig.fir 206131:4]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:19 chipyard.TestHarness.TinyRocketConfig.fir 206132:4 Reg.scala 16:23 chipyard.TestHarness.TinyRocketConfig.fir 206133:6 Reg.scala 15:16 chipyard.TestHarness.TinyRocketConfig.fir 206131:4]
  wire  bundleOut_0_a_bits_source_hi_lo = ~_GEN_5; // @[Fragmenter.scala 297:23 chipyard.TestHarness.TinyRocketConfig.fir 206136:4]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 Fragmenter.scala 303:15 chipyard.TestHarness.TinyRocketConfig.fir 206145:4]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 206137:4]
  wire  _repeater_io_repeat_T = ~aHasData; // @[Fragmenter.scala 302:31 chipyard.TestHarness.TinyRocketConfig.fir 206141:4]
  wire  _repeater_io_repeat_T_1 = new_gennum != 4'h0; // @[Fragmenter.scala 302:53 chipyard.TestHarness.TinyRocketConfig.fir 206142:4]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 2'h0}; // @[Fragmenter.scala 304:65 chipyard.TestHarness.TinyRocketConfig.fir 206146:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90 chipyard.TestHarness.TinyRocketConfig.fir 206147:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88 chipyard.TestHarness.TinyRocketConfig.fir 206148:4]
  wire [5:0] _GEN_10 = {{4'd0}, aFragOH1}; // @[Fragmenter.scala 304:100 chipyard.TestHarness.TinyRocketConfig.fir 206149:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10; // @[Fragmenter.scala 304:100 chipyard.TestHarness.TinyRocketConfig.fir 206149:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h3; // @[Fragmenter.scala 304:111 chipyard.TestHarness.TinyRocketConfig.fir 206150:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51 chipyard.TestHarness.TinyRocketConfig.fir 206151:4]
  wire [28:0] _GEN_11 = {{23'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49 chipyard.TestHarness.TinyRocketConfig.fir 206152:4]
  wire [2:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,bundleOut_0_a_bits_source_hi_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 206154:4]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17 chipyard.TestHarness.TinyRocketConfig.fir 206158:4]
  wire  _T_11 = _T_9 | _repeater_io_repeat_T; // @[Fragmenter.scala 309:35 chipyard.TestHarness.TinyRocketConfig.fir 206160:4]
  wire  _T_13 = _T_11 | reset; // @[Fragmenter.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206162:4]
  wire  _T_14 = ~_T_13; // @[Fragmenter.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206163:4]
  wire  _T_16 = repeater_io_deq_bits_mask == 4'hf; // @[Fragmenter.scala 312:53 chipyard.TestHarness.TinyRocketConfig.fir 206170:4]
  wire  _T_17 = _T_9 | _T_16; // @[Fragmenter.scala 312:35 chipyard.TestHarness.TinyRocketConfig.fir 206171:4]
  wire  _T_19 = _T_17 | reset; // @[Fragmenter.scala 312:16 chipyard.TestHarness.TinyRocketConfig.fir 206173:4]
  wire  _T_20 = ~_T_19; // @[Fragmenter.scala 312:16 chipyard.TestHarness.TinyRocketConfig.fir 206174:4]
  TLMonitor_44_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 205975:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Repeater_7_inTestHarness repeater ( // @[Fragmenter.scala 262:30 chipyard.TestHarness.TinyRocketConfig.fir 206077:4]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_opcode(repeater_io_enq_bits_opcode),
    .io_enq_bits_param(repeater_io_enq_bits_param),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_opcode(repeater_io_deq_bits_opcode),
    .io_deq_bits_param(repeater_io_deq_bits_param),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 Fragmenter.scala 263:25 chipyard.TestHarness.TinyRocketConfig.fir 206081:4]
  assign auto_in_d_valid = auto_out_d_valid & _bundleIn_0_d_valid_T; // @[Fragmenter.scala 224:36 chipyard.TestHarness.TinyRocketConfig.fir 206070:4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32 chipyard.TestHarness.TinyRocketConfig.fir 206075:4]
  assign auto_in_d_bits_source = auto_out_d_bits_source[6:5]; // @[Fragmenter.scala 226:47 chipyard.TestHarness.TinyRocketConfig.fir 206073:4]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 Fragmenter.scala 303:15 chipyard.TestHarness.TinyRocketConfig.fir 206145:4]
  assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 Fragmenter.scala 303:15 chipyard.TestHarness.TinyRocketConfig.fir 206145:4]
  assign auto_out_a_bits_param = repeater_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 Fragmenter.scala 303:15 chipyard.TestHarness.TinyRocketConfig.fir 206145:4]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 Fragmenter.scala 306:25 chipyard.TestHarness.TinyRocketConfig.fir 206157:4]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 206155:4]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11; // @[Fragmenter.scala 304:49 chipyard.TestHarness.TinyRocketConfig.fir 206152:4]
  assign auto_out_a_bits_mask = repeater_io_full ? 4'hf : auto_in_a_bits_mask; // @[Fragmenter.scala 313:31 chipyard.TestHarness.TinyRocketConfig.fir 206179:4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 Fragmenter.scala 303:15 chipyard.TestHarness.TinyRocketConfig.fir 206145:4]
  assign auto_out_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35 chipyard.TestHarness.TinyRocketConfig.fir 206067:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 205976:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 205977:4]
  assign monitor_io_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 Fragmenter.scala 263:25 chipyard.TestHarness.TinyRocketConfig.fir 206081:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign monitor_io_in_d_valid = auto_out_d_valid & _bundleIn_0_d_valid_T; // @[Fragmenter.scala 224:36 chipyard.TestHarness.TinyRocketConfig.fir 206070:4]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign monitor_io_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32 chipyard.TestHarness.TinyRocketConfig.fir 206075:4]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source[6:5]; // @[Fragmenter.scala 226:47 chipyard.TestHarness.TinyRocketConfig.fir 206073:4]
  assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  assign repeater_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 206079:4]
  assign repeater_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 206080:4]
  assign repeater_io_repeat = _repeater_io_repeat_T & _repeater_io_repeat_T_1; // @[Fragmenter.scala 302:41 chipyard.TestHarness.TinyRocketConfig.fir 206143:4]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign repeater_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 205973:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206001:4]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 205998:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 206000:4]
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29 chipyard.TestHarness.TinyRocketConfig.fir 206002:4]
      acknum <= 4'h0; // @[Fragmenter.scala 189:29 chipyard.TestHarness.TinyRocketConfig.fir 206002:4]
    end else if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.TinyRocketConfig.fir 206052:4]
      if (dFirst) begin // @[Fragmenter.scala 209:24 chipyard.TestHarness.TinyRocketConfig.fir 206055:6]
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.TinyRocketConfig.fir 206052:4]
      if (dFirst) begin // @[Fragmenter.scala 210:25 chipyard.TestHarness.TinyRocketConfig.fir 206057:6]
        dOrig <= dFirst_size; // @[Fragmenter.scala 211:19 chipyard.TestHarness.TinyRocketConfig.fir 206058:8]
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30 chipyard.TestHarness.TinyRocketConfig.fir 206004:4]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30 chipyard.TestHarness.TinyRocketConfig.fir 206004:4]
    end else if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.TinyRocketConfig.fir 206052:4]
      if (dFirst) begin // @[Fragmenter.scala 210:25 chipyard.TestHarness.TinyRocketConfig.fir 206057:6]
        dToggle <= auto_out_d_bits_source[4]; // @[Fragmenter.scala 212:21 chipyard.TestHarness.TinyRocketConfig.fir 206060:8]
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29 chipyard.TestHarness.TinyRocketConfig.fir 206115:4]
      gennum <= 4'h0; // @[Fragmenter.scala 291:29 chipyard.TestHarness.TinyRocketConfig.fir 206115:4]
    end else if (_T_8) begin // @[Fragmenter.scala 300:29 chipyard.TestHarness.TinyRocketConfig.fir 206138:4]
      gennum <= new_gennum; // @[Fragmenter.scala 300:38 chipyard.TestHarness.TinyRocketConfig.fir 206139:6]
    end
    if (aFirst) begin // @[Reg.scala 16:19 chipyard.TestHarness.TinyRocketConfig.fir 206132:4]
      aToggle_r <= dToggle; // @[Reg.scala 16:23 chipyard.TestHarness.TinyRocketConfig.fir 206133:6]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:309 assert (!repeater.io.full || !aHasData)\n"
            ); // @[Fragmenter.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206165:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_14) begin
          $fatal; // @[Fragmenter.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 206166:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16 chipyard.TestHarness.TinyRocketConfig.fir 206176:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_20) begin
          $fatal; // @[Fragmenter.scala 312:16 chipyard.TestHarness.TinyRocketConfig.fir 206177:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_45_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 206217:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 206218:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 206219:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input  [3:0]  io_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input  [31:0] io_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input  [3:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input  [3:0]  io_in_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input         io_in_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input         io_in_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 206220:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 208057:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 208364:4]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 206236:6]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 206238:6]
  wire [31:0] _GEN_71 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.TinyRocketConfig.fir 206239:6]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.TinyRocketConfig.fir 206239:6]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24 chipyard.TestHarness.TinyRocketConfig.fir 206240:6]
  wire  mask_sizeOH_shiftAmount = io_in_a_bits_size[0]; // @[OneHot.scala 64:49 chipyard.TestHarness.TinyRocketConfig.fir 206242:6]
  wire [1:0] _mask_sizeOH_T_1 = 2'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.TinyRocketConfig.fir 206243:6]
  wire [1:0] mask_sizeOH = _mask_sizeOH_T_1 | 2'h1; // @[Misc.scala 201:81 chipyard.TestHarness.TinyRocketConfig.fir 206245:6]
  wire  _mask_T = io_in_a_bits_size >= 4'h2; // @[Misc.scala 205:21 chipyard.TestHarness.TinyRocketConfig.fir 206246:6]
  wire  mask_size = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 206247:6]
  wire  mask_bit = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 206248:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 206249:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 206251:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 206252:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 206254:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 206255:6]
  wire  mask_size_1 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.TinyRocketConfig.fir 206256:6]
  wire  mask_bit_1 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.TinyRocketConfig.fir 206257:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.TinyRocketConfig.fir 206258:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 206259:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 206260:6]
  wire  mask_lo_lo = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 206261:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 206262:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 206263:6]
  wire  mask_lo_hi = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 206264:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 206265:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 206266:6]
  wire  mask_hi_lo = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 206267:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.TinyRocketConfig.fir 206268:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.TinyRocketConfig.fir 206269:6]
  wire  mask_hi_hi = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.TinyRocketConfig.fir 206270:6]
  wire [3:0] mask = {mask_hi_hi,mask_hi_lo,mask_lo_hi,mask_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.TinyRocketConfig.fir 206273:6]
  wire [32:0] _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 206277:6]
  wire  _T_15 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.TinyRocketConfig.fir 206289:6]
  wire  _T_17 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42 chipyard.TestHarness.TinyRocketConfig.fir 206292:8]
  wire [32:0] _T_26 = $signed(_T_7) & -33'sh101000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 206301:8]
  wire  _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 206302:8]
  wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 206303:8]
  wire [32:0] _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 206304:8]
  wire [32:0] _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 206306:8]
  wire  _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 206307:8]
  wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 206308:8]
  wire [32:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 206309:8]
  wire [32:0] _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 206311:8]
  wire  _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 206312:8]
  wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 206313:8]
  wire [32:0] _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 206314:8]
  wire [32:0] _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 206316:8]
  wire  _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 206317:8]
  wire [31:0] _T_43 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 206318:8]
  wire [32:0] _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 206319:8]
  wire [32:0] _T_46 = $signed(_T_44) & -33'sh4000000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 206321:8]
  wire  _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 206322:8]
  wire [31:0] _T_48 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 206323:8]
  wire [32:0] _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 206324:8]
  wire [32:0] _T_51 = $signed(_T_49) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 206326:8]
  wire  _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 206327:8]
  wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h54000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 206328:8]
  wire [32:0] _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 206329:8]
  wire [32:0] _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 206331:8]
  wire  _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 206332:8]
  wire [31:0] _T_58 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31 chipyard.TestHarness.TinyRocketConfig.fir 206333:8]
  wire [32:0] _T_59 = {1'b0,$signed(_T_58)}; // @[Parameters.scala 137:49 chipyard.TestHarness.TinyRocketConfig.fir 206334:8]
  wire [32:0] _T_61 = $signed(_T_59) & -33'sh4000; // @[Parameters.scala 137:52 chipyard.TestHarness.TinyRocketConfig.fir 206336:8]
  wire  _T_62 = $signed(_T_61) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.TinyRocketConfig.fir 206337:8]
  wire  _T_63 = _T_27 | _T_32; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206338:8]
  wire  _T_75 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206350:8]
  wire  _T_138 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206425:8]
  wire  _T_139 = ~_T_138; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206426:8]
  wire  _T_141 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206432:8]
  wire  _T_142 = ~_T_141; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206433:8]
  wire [3:0] _T_147 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.TinyRocketConfig.fir 206446:8]
  wire  _T_148 = _T_147 == 4'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.TinyRocketConfig.fir 206447:8]
  wire  _T_150 = _T_148 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206449:8]
  wire  _T_151 = ~_T_150; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206450:8]
  wire  _T_156 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.TinyRocketConfig.fir 206464:6]
  wire  _T_301 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.TinyRocketConfig.fir 206647:6]
  wire  _T_309 = _T_17 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206656:8]
  wire  _T_310 = ~_T_309; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206657:8]
  wire  _T_320 = _T_17 & _T_32; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 206671:8]
  wire  _T_322 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.TinyRocketConfig.fir 206673:8]
  wire  _T_360 = _T_27 | _T_37; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206711:8]
  wire  _T_361 = _T_360 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206712:8]
  wire  _T_362 = _T_361 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206713:8]
  wire  _T_363 = _T_362 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206714:8]
  wire  _T_364 = _T_363 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206715:8]
  wire  _T_365 = _T_364 | _T_62; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206716:8]
  wire  _T_366 = _T_322 & _T_365; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 206717:8]
  wire  _T_368 = _T_320 | _T_366; // @[Parameters.scala 672:30 chipyard.TestHarness.TinyRocketConfig.fir 206719:8]
  wire  _T_370 = _T_368 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206721:8]
  wire  _T_371 = ~_T_370; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206722:8]
  wire  _T_382 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.TinyRocketConfig.fir 206749:8]
  wire  _T_384 = _T_382 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206751:8]
  wire  _T_385 = ~_T_384; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206752:8]
  wire  _T_390 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.TinyRocketConfig.fir 206766:6]
  wire  _T_441 = _T_27 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206818:8]
  wire  _T_442 = _T_441 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206819:8]
  wire  _T_443 = _T_442 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206820:8]
  wire  _T_444 = _T_443 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206821:8]
  wire  _T_445 = _T_444 | _T_62; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 206822:8]
  wire  _T_446 = _T_322 & _T_445; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 206823:8]
  wire  _T_455 = _T_320 | _T_446; // @[Parameters.scala 672:30 chipyard.TestHarness.TinyRocketConfig.fir 206832:8]
  wire  _T_457 = _T_17 & _T_455; // @[Monitor.scala 115:71 chipyard.TestHarness.TinyRocketConfig.fir 206834:8]
  wire  _T_459 = _T_457 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206836:8]
  wire  _T_460 = ~_T_459; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206837:8]
  wire  _T_475 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.TinyRocketConfig.fir 206873:6]
  wire [3:0] _T_556 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.TinyRocketConfig.fir 206971:8]
  wire [3:0] _T_557 = io_in_a_bits_mask & _T_556; // @[Monitor.scala 127:31 chipyard.TestHarness.TinyRocketConfig.fir 206972:8]
  wire  _T_558 = _T_557 == 4'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.TinyRocketConfig.fir 206973:8]
  wire  _T_560 = _T_558 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206975:8]
  wire  _T_561 = ~_T_560; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206976:8]
  wire  _T_562 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.TinyRocketConfig.fir 206982:6]
  wire  _T_570 = io_in_a_bits_size <= 4'h2; // @[Parameters.scala 92:42 chipyard.TestHarness.TinyRocketConfig.fir 206991:8]
  wire  _T_609 = _T_63 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 207030:8]
  wire  _T_610 = _T_609 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 207031:8]
  wire  _T_611 = _T_610 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 207032:8]
  wire  _T_612 = _T_611 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 207033:8]
  wire  _T_613 = _T_612 | _T_62; // @[Parameters.scala 671:42 chipyard.TestHarness.TinyRocketConfig.fir 207034:8]
  wire  _T_614 = _T_570 & _T_613; // @[Parameters.scala 670:56 chipyard.TestHarness.TinyRocketConfig.fir 207035:8]
  wire  _T_624 = _T_17 & _T_614; // @[Monitor.scala 131:74 chipyard.TestHarness.TinyRocketConfig.fir 207045:8]
  wire  _T_626 = _T_624 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207047:8]
  wire  _T_627 = ~_T_626; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207048:8]
  wire  _T_642 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.TinyRocketConfig.fir 207084:6]
  wire  _T_722 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.TinyRocketConfig.fir 207186:6]
  wire  _T_784 = _T_17 & _T_320; // @[Monitor.scala 147:68 chipyard.TestHarness.TinyRocketConfig.fir 207249:8]
  wire  _T_786 = _T_784 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207251:8]
  wire  _T_787 = ~_T_786; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207252:8]
  wire  _T_806 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.TinyRocketConfig.fir 207298:6]
  wire  _T_808 = _T_806 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207300:6]
  wire  _T_809 = ~_T_808; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207301:6]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.TinyRocketConfig.fir 207306:6]
  wire  _T_810 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.TinyRocketConfig.fir 207311:6]
  wire  _T_812 = _source_ok_T_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207314:8]
  wire  _T_813 = ~_T_812; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207315:8]
  wire  _T_814 = io_in_d_bits_size >= 4'h2; // @[Monitor.scala 312:27 chipyard.TestHarness.TinyRocketConfig.fir 207320:8]
  wire  _T_816 = _T_814 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207322:8]
  wire  _T_817 = ~_T_816; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207323:8]
  wire  _T_818 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.TinyRocketConfig.fir 207328:8]
  wire  _T_820 = _T_818 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207330:8]
  wire  _T_821 = ~_T_820; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207331:8]
  wire  _T_822 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.TinyRocketConfig.fir 207336:8]
  wire  _T_824 = _T_822 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207338:8]
  wire  _T_825 = ~_T_824; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207339:8]
  wire  _T_826 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.TinyRocketConfig.fir 207344:8]
  wire  _T_828 = _T_826 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207346:8]
  wire  _T_829 = ~_T_828; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207347:8]
  wire  _T_830 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.TinyRocketConfig.fir 207353:6]
  wire  _T_841 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.TinyRocketConfig.fir 207377:8]
  wire  _T_843 = _T_841 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207379:8]
  wire  _T_844 = ~_T_843; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207380:8]
  wire  _T_845 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.TinyRocketConfig.fir 207385:8]
  wire  _T_847 = _T_845 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207387:8]
  wire  _T_848 = ~_T_847; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207388:8]
  wire  _T_858 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.TinyRocketConfig.fir 207411:6]
  wire  _T_878 = _T_826 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.TinyRocketConfig.fir 207452:8]
  wire  _T_880 = _T_878 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207454:8]
  wire  _T_881 = ~_T_880; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207455:8]
  wire  _T_887 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.TinyRocketConfig.fir 207470:6]
  wire  _T_904 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.TinyRocketConfig.fir 207505:6]
  wire  _T_922 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.TinyRocketConfig.fir 207541:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 207607:4]
  wire [9:0] a_first_beats1_decode = is_aligned_mask[11:2]; // @[Edges.scala 219:59 chipyard.TestHarness.TinyRocketConfig.fir 207612:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.TinyRocketConfig.fir 207614:4]
  reg [9:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207616:4]
  wire [9:0] a_first_counter1 = a_first_counter - 10'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 207618:4]
  wire  a_first = a_first_counter == 10'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 207619:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.TinyRocketConfig.fir 207630:4]
  reg [3:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.TinyRocketConfig.fir 207632:4]
  reg [31:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.TinyRocketConfig.fir 207634:4]
  wire  _T_951 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.TinyRocketConfig.fir 207635:4]
  wire  _T_952 = io_in_a_valid & _T_951; // @[Monitor.scala 389:19 chipyard.TestHarness.TinyRocketConfig.fir 207636:4]
  wire  _T_953 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.TinyRocketConfig.fir 207638:6]
  wire  _T_955 = _T_953 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207640:6]
  wire  _T_956 = ~_T_955; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207641:6]
  wire  _T_961 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.TinyRocketConfig.fir 207654:6]
  wire  _T_963 = _T_961 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207656:6]
  wire  _T_964 = ~_T_963; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207657:6]
  wire  _T_969 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.TinyRocketConfig.fir 207670:6]
  wire  _T_971 = _T_969 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207672:6]
  wire  _T_972 = ~_T_971; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207673:6]
  wire  _T_974 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.TinyRocketConfig.fir 207680:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 207688:4]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.TinyRocketConfig.fir 207690:4]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.TinyRocketConfig.fir 207692:4]
  wire [9:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:2]; // @[Edges.scala 219:59 chipyard.TestHarness.TinyRocketConfig.fir 207693:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.TinyRocketConfig.fir 207694:4]
  reg [9:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207696:4]
  wire [9:0] d_first_counter1 = d_first_counter - 10'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 207698:4]
  wire  d_first = d_first_counter == 10'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 207699:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.TinyRocketConfig.fir 207710:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.TinyRocketConfig.fir 207711:4]
  reg [3:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.TinyRocketConfig.fir 207712:4]
  reg  source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.TinyRocketConfig.fir 207713:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.TinyRocketConfig.fir 207714:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.TinyRocketConfig.fir 207715:4]
  wire  _T_975 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.TinyRocketConfig.fir 207716:4]
  wire  _T_976 = io_in_d_valid & _T_975; // @[Monitor.scala 541:19 chipyard.TestHarness.TinyRocketConfig.fir 207717:4]
  wire  _T_977 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.TinyRocketConfig.fir 207719:6]
  wire  _T_979 = _T_977 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207721:6]
  wire  _T_980 = ~_T_979; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207722:6]
  wire  _T_981 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.TinyRocketConfig.fir 207727:6]
  wire  _T_983 = _T_981 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207729:6]
  wire  _T_984 = ~_T_983; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207730:6]
  wire  _T_985 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.TinyRocketConfig.fir 207735:6]
  wire  _T_987 = _T_985 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207737:6]
  wire  _T_988 = ~_T_987; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207738:6]
  wire  _T_989 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.TinyRocketConfig.fir 207743:6]
  wire  _T_991 = _T_989 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207745:6]
  wire  _T_992 = ~_T_991; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207746:6]
  wire  _T_993 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.TinyRocketConfig.fir 207751:6]
  wire  _T_995 = _T_993 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207753:6]
  wire  _T_996 = ~_T_995; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207754:6]
  wire  _T_997 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.TinyRocketConfig.fir 207759:6]
  wire  _T_999 = _T_997 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207761:6]
  wire  _T_1000 = ~_T_999; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207762:6]
  wire  _T_1002 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.TinyRocketConfig.fir 207769:4]
  reg  inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 207778:4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 207779:4]
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 207780:4]
  reg [9:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207790:4]
  wire [9:0] a_first_counter1_1 = a_first_counter_1 - 10'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 207792:4]
  wire  a_first_1 = a_first_counter_1 == 10'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 207793:4]
  reg [9:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207812:4]
  wire [9:0] d_first_counter1_1 = d_first_counter_1 - 10'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 207814:4]
  wire  d_first_1 = d_first_counter_1 == 10'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 207815:4]
  wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.TinyRocketConfig.fir 207836:4]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.TinyRocketConfig.fir 207836:4]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.TinyRocketConfig.fir 207837:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.TinyRocketConfig.fir 207841:4]
  wire [15:0] _GEN_73 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.TinyRocketConfig.fir 207842:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.TinyRocketConfig.fir 207842:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.TinyRocketConfig.fir 207843:4]
  wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65 chipyard.TestHarness.TinyRocketConfig.fir 207847:4]
  wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.TinyRocketConfig.fir 207848:4]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.TinyRocketConfig.fir 207852:4]
  wire [15:0] _GEN_75 = {{8'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.TinyRocketConfig.fir 207853:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.TinyRocketConfig.fir 207853:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.TinyRocketConfig.fir 207854:4]
  wire  _T_1003 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.TinyRocketConfig.fir 207878:4]
  wire [1:0] _GEN_15 = _T_1003 ? 2'h1 : 2'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.TinyRocketConfig.fir 207880:4 Monitor.scala 649:22 chipyard.TestHarness.TinyRocketConfig.fir 207882:6 chipyard.TestHarness.TinyRocketConfig.fir 207829:4]
  wire  _T_1006 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.TinyRocketConfig.fir 207885:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.TinyRocketConfig.fir 207890:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.TinyRocketConfig.fir 207891:6]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.TinyRocketConfig.fir 207893:6]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.TinyRocketConfig.fir 207894:6]
  wire [3:0] a_opcodes_set_interm = _T_1006 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 207887:4 Monitor.scala 654:28 chipyard.TestHarness.TinyRocketConfig.fir 207892:6 chipyard.TestHarness.TinyRocketConfig.fir 207875:4]
  wire [18:0] _a_opcodes_set_T_1 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.TinyRocketConfig.fir 207897:6]
  wire [4:0] a_sizes_set_interm = _T_1006 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 207887:4 Monitor.scala 655:28 chipyard.TestHarness.TinyRocketConfig.fir 207895:6 chipyard.TestHarness.TinyRocketConfig.fir 207877:4]
  wire [19:0] _a_sizes_set_T_1 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.TinyRocketConfig.fir 207900:6]
  wire  _T_1010 = ~inflight; // @[Monitor.scala 658:17 chipyard.TestHarness.TinyRocketConfig.fir 207904:6]
  wire  _T_1012 = _T_1010 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207906:6]
  wire  _T_1013 = ~_T_1012; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207907:6]
  wire [1:0] _GEN_16 = _T_1006 ? 2'h1 : 2'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 207887:4 Monitor.scala 653:28 chipyard.TestHarness.TinyRocketConfig.fir 207889:6 chipyard.TestHarness.TinyRocketConfig.fir 207827:4]
  wire [18:0] _GEN_19 = _T_1006 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 207887:4 Monitor.scala 656:28 chipyard.TestHarness.TinyRocketConfig.fir 207898:6 chipyard.TestHarness.TinyRocketConfig.fir 207831:4]
  wire [19:0] _GEN_20 = _T_1006 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.TinyRocketConfig.fir 207887:4 Monitor.scala 657:28 chipyard.TestHarness.TinyRocketConfig.fir 207901:6 chipyard.TestHarness.TinyRocketConfig.fir 207833:4]
  wire  _T_1014 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.TinyRocketConfig.fir 207922:4]
  wire  _T_1016 = ~_T_810; // @[Monitor.scala 671:74 chipyard.TestHarness.TinyRocketConfig.fir 207924:4]
  wire  _T_1017 = _T_1014 & _T_1016; // @[Monitor.scala 671:71 chipyard.TestHarness.TinyRocketConfig.fir 207925:4]
  wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.TinyRocketConfig.fir 207927:6]
  wire [1:0] _GEN_21 = _T_1017 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.TinyRocketConfig.fir 207926:4 Monitor.scala 672:22 chipyard.TestHarness.TinyRocketConfig.fir 207928:6 chipyard.TestHarness.TinyRocketConfig.fir 207916:4]
  wire  _T_1019 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.TinyRocketConfig.fir 207931:4]
  wire  _T_1022 = _T_1019 & _T_1016; // @[Monitor.scala 675:72 chipyard.TestHarness.TinyRocketConfig.fir 207934:4]
  wire [30:0] _GEN_78 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.TinyRocketConfig.fir 207943:6]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_78 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.TinyRocketConfig.fir 207943:6]
  wire [30:0] _GEN_79 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74 chipyard.TestHarness.TinyRocketConfig.fir 207950:6]
  wire [30:0] _d_sizes_clr_T_5 = _GEN_79 << _a_size_lookup_T; // @[Monitor.scala 678:74 chipyard.TestHarness.TinyRocketConfig.fir 207950:6]
  wire [1:0] _GEN_22 = _T_1022 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 207935:4 Monitor.scala 676:21 chipyard.TestHarness.TinyRocketConfig.fir 207937:6 chipyard.TestHarness.TinyRocketConfig.fir 207914:4]
  wire [30:0] _GEN_23 = _T_1022 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 207935:4 Monitor.scala 677:21 chipyard.TestHarness.TinyRocketConfig.fir 207944:6 chipyard.TestHarness.TinyRocketConfig.fir 207918:4]
  wire [30:0] _GEN_24 = _T_1022 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.TinyRocketConfig.fir 207935:4 Monitor.scala 678:21 chipyard.TestHarness.TinyRocketConfig.fir 207951:6 chipyard.TestHarness.TinyRocketConfig.fir 207920:4]
  wire  same_cycle_resp = _T_1003 & _source_ok_T_1; // @[Monitor.scala 681:88 chipyard.TestHarness.TinyRocketConfig.fir 207961:6]
  wire  _T_1027 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.TinyRocketConfig.fir 207962:6]
  wire  _T_1029 = _T_1027 | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.TinyRocketConfig.fir 207964:6]
  wire  _T_1031 = _T_1029 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207966:6]
  wire  _T_1032 = ~_T_1031; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207967:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8 Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8]
  wire  _T_1033 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.TinyRocketConfig.fir 207973:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 207974:8 Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 207974:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 207974:8 Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 207974:8]
  wire  _T_1034 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.TinyRocketConfig.fir 207974:8]
  wire  _T_1035 = _T_1033 | _T_1034; // @[Monitor.scala 685:77 chipyard.TestHarness.TinyRocketConfig.fir 207975:8]
  wire  _T_1037 = _T_1035 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207977:8]
  wire  _T_1038 = ~_T_1037; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207978:8]
  wire  _T_1039 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.TinyRocketConfig.fir 207983:8]
  wire  _T_1041 = _T_1039 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207985:8]
  wire  _T_1042 = ~_T_1041; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207986:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 207834:4 Monitor.scala 634:21 chipyard.TestHarness.TinyRocketConfig.fir 207844:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8 Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8]
  wire  _T_1044 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.TinyRocketConfig.fir 207994:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 207996:8 Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 207996:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 207996:8 Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 207996:8]
  wire  _T_1046 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.TinyRocketConfig.fir 207996:8]
  wire  _T_1047 = _T_1044 | _T_1046; // @[Monitor.scala 689:72 chipyard.TestHarness.TinyRocketConfig.fir 207997:8]
  wire  _T_1049 = _T_1047 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207999:8]
  wire  _T_1050 = ~_T_1049; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208000:8]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 207845:4 Monitor.scala 638:19 chipyard.TestHarness.TinyRocketConfig.fir 207855:4]
  wire [7:0] _GEN_80 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.TinyRocketConfig.fir 208005:8]
  wire  _T_1051 = _GEN_80 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.TinyRocketConfig.fir 208005:8]
  wire  _T_1053 = _T_1051 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208007:8]
  wire  _T_1054 = ~_T_1053; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208008:8]
  wire  _T_1056 = _T_1014 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.TinyRocketConfig.fir 208016:4]
  wire  _T_1057 = _T_1056 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.TinyRocketConfig.fir 208017:4]
  wire  _T_1059 = _T_1057 & _source_ok_T_1; // @[Monitor.scala 694:65 chipyard.TestHarness.TinyRocketConfig.fir 208019:4]
  wire  _T_1061 = _T_1059 & _T_1016; // @[Monitor.scala 694:116 chipyard.TestHarness.TinyRocketConfig.fir 208021:4]
  wire  _T_1062 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.TinyRocketConfig.fir 208023:6]
  wire  _T_1063 = _T_1062 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.TinyRocketConfig.fir 208024:6]
  wire  _T_1065 = _T_1063 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208026:6]
  wire  _T_1066 = ~_T_1065; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208027:6]
  wire  a_set_wo_ready = _GEN_15[0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 207828:4]
  wire  d_clr_wo_ready = _GEN_21[0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 207915:4]
  wire  _T_1067 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.TinyRocketConfig.fir 208033:4]
  wire  _T_1068 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.TinyRocketConfig.fir 208034:4]
  wire  _T_1069 = ~_T_1068; // @[Monitor.scala 699:51 chipyard.TestHarness.TinyRocketConfig.fir 208035:4]
  wire  _T_1070 = _T_1067 | _T_1069; // @[Monitor.scala 699:48 chipyard.TestHarness.TinyRocketConfig.fir 208036:4]
  wire  _T_1072 = _T_1070 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208038:4]
  wire  _T_1073 = ~_T_1072; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208039:4]
  wire  a_set = _GEN_16[0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 207826:4]
  wire  _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.TinyRocketConfig.fir 208044:4]
  wire  d_clr = _GEN_22[0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 207913:4]
  wire  _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.TinyRocketConfig.fir 208045:4]
  wire  _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.TinyRocketConfig.fir 208046:4]
  wire [3:0] a_opcodes_set = _GEN_19[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 207830:4]
  wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.TinyRocketConfig.fir 208048:4]
  wire [3:0] d_opcodes_clr = _GEN_23[3:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 207917:4]
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.TinyRocketConfig.fir 208049:4]
  wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.TinyRocketConfig.fir 208050:4]
  wire [7:0] a_sizes_set = _GEN_20[7:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 207832:4]
  wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.TinyRocketConfig.fir 208052:4]
  wire [7:0] d_sizes_clr = _GEN_24[7:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 207919:4]
  wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56 chipyard.TestHarness.TinyRocketConfig.fir 208053:4]
  wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.TinyRocketConfig.fir 208054:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 208056:4]
  wire  _T_1074 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.TinyRocketConfig.fir 208059:4]
  wire  _T_1075 = ~_T_1074; // @[Monitor.scala 709:16 chipyard.TestHarness.TinyRocketConfig.fir 208060:4]
  wire  _T_1076 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.TinyRocketConfig.fir 208061:4]
  wire  _T_1077 = _T_1075 | _T_1076; // @[Monitor.scala 709:30 chipyard.TestHarness.TinyRocketConfig.fir 208062:4]
  wire  _T_1078 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.TinyRocketConfig.fir 208063:4]
  wire  _T_1079 = _T_1077 | _T_1078; // @[Monitor.scala 709:47 chipyard.TestHarness.TinyRocketConfig.fir 208064:4]
  wire  _T_1081 = _T_1079 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 208066:4]
  wire  _T_1082 = ~_T_1081; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 208067:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.TinyRocketConfig.fir 208073:4]
  wire  _T_1085 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.TinyRocketConfig.fir 208077:4]
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 208083:4]
  reg [9:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 208118:4]
  wire [9:0] d_first_counter1_2 = d_first_counter_2 - 10'h1; // @[Edges.scala 229:28 chipyard.TestHarness.TinyRocketConfig.fir 208120:4]
  wire  d_first_2 = d_first_counter_2 == 10'h0; // @[Edges.scala 230:25 chipyard.TestHarness.TinyRocketConfig.fir 208121:4]
  wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.TinyRocketConfig.fir 208154:4]
  wire [15:0] _GEN_84 = {{8'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.TinyRocketConfig.fir 208159:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_84 & _a_size_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.TinyRocketConfig.fir 208159:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.TinyRocketConfig.fir 208160:4]
  wire  _T_1103 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.TinyRocketConfig.fir 208238:4]
  wire  _T_1105 = _T_1103 & _T_810; // @[Monitor.scala 779:71 chipyard.TestHarness.TinyRocketConfig.fir 208240:4]
  wire  _T_1107 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.TinyRocketConfig.fir 208246:4]
  wire  _T_1109 = _T_1107 & _T_810; // @[Monitor.scala 783:72 chipyard.TestHarness.TinyRocketConfig.fir 208248:4]
  wire [30:0] _GEN_69 = _T_1109 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.TinyRocketConfig.fir 208249:4 Monitor.scala 786:21 chipyard.TestHarness.TinyRocketConfig.fir 208265:6 chipyard.TestHarness.TinyRocketConfig.fir 208236:4]
  wire  _T_1113 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.TinyRocketConfig.fir 208284:6]
  wire  _T_1117 = _T_1113 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208288:6]
  wire  _T_1118 = ~_T_1117; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208289:6]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 208142:4 Monitor.scala 747:21 chipyard.TestHarness.TinyRocketConfig.fir 208161:4]
  wire  _T_1123 = _GEN_80 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.TinyRocketConfig.fir 208307:8]
  wire  _T_1125 = _T_1123 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208309:8]
  wire  _T_1126 = ~_T_1125; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208310:8]
  wire [7:0] d_sizes_clr_1 = _GEN_69[7:0]; // @[chipyard.TestHarness.TinyRocketConfig.fir 208235:4]
  wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58 chipyard.TestHarness.TinyRocketConfig.fir 208360:4]
  wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.TinyRocketConfig.fir 208361:4]
  wire  _GEN_90 = io_in_a_valid & _T_15; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206352:10]
  wire  _GEN_100 = io_in_a_valid & _T_156; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206527:10]
  wire  _GEN_112 = io_in_a_valid & _T_301; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206659:10]
  wire  _GEN_120 = io_in_a_valid & _T_390; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206839:10]
  wire  _GEN_126 = io_in_a_valid & _T_475; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206946:10]
  wire  _GEN_132 = io_in_a_valid & _T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207050:10]
  wire  _GEN_138 = io_in_a_valid & _T_642; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207152:10]
  wire  _GEN_144 = io_in_a_valid & _T_722; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207254:10]
  wire  _GEN_150 = io_in_d_valid & _T_810; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207317:10]
  wire  _GEN_160 = io_in_d_valid & _T_830; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207359:10]
  wire  _GEN_172 = io_in_d_valid & _T_858; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207417:10]
  wire  _GEN_184 = io_in_d_valid & _T_887; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207476:10]
  wire  _GEN_190 = io_in_d_valid & _T_904; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207511:10]
  wire  _GEN_196 = io_in_d_valid & _T_922; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207547:10]
  wire  _GEN_202 = _T_1017 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207980:10]
  wire  _GEN_207 = _T_1017 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208002:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 208057:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 208364:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207616:4]
      a_first_counter <= 10'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207616:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 207626:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 207627:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 207615:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 10'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_974) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 207681:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.TinyRocketConfig.fir 207682:6]
    end
    if (_T_974) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 207681:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.TinyRocketConfig.fir 207684:6]
    end
    if (_T_974) begin // @[Monitor.scala 396:32 chipyard.TestHarness.TinyRocketConfig.fir 207681:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.TinyRocketConfig.fir 207686:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207696:4]
      d_first_counter <= 10'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207696:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 207706:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 207707:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 207695:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 10'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 207770:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.TinyRocketConfig.fir 207771:6]
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 207770:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.TinyRocketConfig.fir 207772:6]
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 207770:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.TinyRocketConfig.fir 207773:6]
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 207770:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.TinyRocketConfig.fir 207774:6]
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 207770:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.TinyRocketConfig.fir 207775:6]
    end
    if (_T_1002) begin // @[Monitor.scala 549:32 chipyard.TestHarness.TinyRocketConfig.fir 207770:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.TinyRocketConfig.fir 207776:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 207778:4]
      inflight <= 1'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.TinyRocketConfig.fir 207778:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.TinyRocketConfig.fir 208047:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 207779:4]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.TinyRocketConfig.fir 207779:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.TinyRocketConfig.fir 208051:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 207780:4]
      inflight_sizes <= 8'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.TinyRocketConfig.fir 207780:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.TinyRocketConfig.fir 208055:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207790:4]
      a_first_counter_1 <= 10'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207790:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 207800:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 207801:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 207615:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 10'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207812:4]
      d_first_counter_1 <= 10'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 207812:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 207822:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 207823:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 207695:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 10'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 208056:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.TinyRocketConfig.fir 208056:4]
    end else if (_T_1085) begin // @[Monitor.scala 712:47 chipyard.TestHarness.TinyRocketConfig.fir 208078:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.TinyRocketConfig.fir 208079:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.TinyRocketConfig.fir 208074:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 208083:4]
      inflight_sizes_1 <= 8'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.TinyRocketConfig.fir 208083:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.TinyRocketConfig.fir 208362:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 208118:4]
      d_first_counter_2 <= 10'h0; // @[Edges.scala 228:27 chipyard.TestHarness.TinyRocketConfig.fir 208118:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.TinyRocketConfig.fir 208128:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.TinyRocketConfig.fir 208129:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.TinyRocketConfig.fir 207695:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 10'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_15 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206352:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_75) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206353:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206413:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_75) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206414:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_139) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206428:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_139) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206429:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206435:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206436:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_151) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206452:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_151) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206453:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_156 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206527:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_75) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206528:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206588:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_75) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206589:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_139) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206603:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_139) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206604:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206610:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206611:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206626:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_75) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206627:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_151) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206635:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_151) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206636:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_301 & _T_310) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206659:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_310) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206660:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_371) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206724:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_371) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206725:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206738:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206739:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_385) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206754:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_385) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206755:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_390 & _T_460) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206839:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_460) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206840:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_120 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206853:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206854:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_120 & _T_385) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206869:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_385) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206870:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_475 & _T_460) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206946:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_460) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206947:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_126 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206960:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206961:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_126 & _T_561) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206978:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_561) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 206979:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_562 & _T_627) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207050:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_627) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207051:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207064:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207065:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_385) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207080:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_385) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207081:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_642 & _T_627) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207152:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_627) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207153:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207166:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207167:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_385) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207182:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_385) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207183:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_722 & _T_787) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207254:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_787) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207255:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_142) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207268:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_142) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207269:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_385) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207284:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_385) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207285:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_809) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207303:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_809) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207304:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_810 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207317:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207318:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_817) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207325:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_817) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207326:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_821) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207333:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_821) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207334:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_825) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207341:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_825) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207342:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_829) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207349:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_829) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207350:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_830 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207359:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207360:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207366:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_75) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207367:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_817) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207374:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_817) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207375:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_844) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207382:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_844) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207383:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_848) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207390:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_848) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207391:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_825) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207398:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_825) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207399:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_858 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207417:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207418:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & _T_75) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207424:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & _T_75) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207425:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & _T_817) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207432:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & _T_817) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207433:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & _T_844) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207440:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & _T_844) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207441:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & _T_848) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207448:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & _T_848) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207449:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & _T_881) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207457:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_172 & _T_881) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207458:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_887 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207476:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_184 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207477:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_184 & _T_821) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207484:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_184 & _T_821) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207485:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_184 & _T_825) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207492:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_184 & _T_825) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207493:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_904 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207511:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_190 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207512:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_190 & _T_821) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207519:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_190 & _T_821) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207520:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_190 & _T_881) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207528:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_190 & _T_881) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207529:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_922 & _T_813) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207547:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_196 & _T_813) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207548:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_196 & _T_821) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207555:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_196 & _T_821) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207556:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_196 & _T_825) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207563:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_196 & _T_825) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207564:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_952 & _T_956) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207643:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_952 & _T_956) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207644:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_952 & _T_964) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207659:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_952 & _T_964) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207660:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_952 & _T_972) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207675:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_952 & _T_972) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207676:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_980) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207724:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_980) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207725:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_984) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207732:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_984) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207733:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_988) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207740:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_988) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207741:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_992) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207748:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_992) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207749:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_996) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207756:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_996) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207757:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_976 & _T_1000) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207764:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_976 & _T_1000) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207765:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1006 & _T_1013) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207909:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1006 & _T_1013) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 207910:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1017 & _T_1032) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207969:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1017 & _T_1032) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207970:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1017 & same_cycle_resp & _T_1038) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207980:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_1038) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207981:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_1042) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207988:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_1042) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 207989:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1017 & ~same_cycle_resp & _T_1050) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208002:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_207 & _T_1050) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208003:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_207 & _T_1054) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208010:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_207 & _T_1054) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208011:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1061 & _T_1066) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208029:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1061 & _T_1066) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208030:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1073) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 8 (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208041:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1073) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208042:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1082) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 208069:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1082) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.TinyRocketConfig.fir 208070:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1105 & _T_1118) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208291:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1105 & _T_1118) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208292:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1105 & _T_1126) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208312:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1105 & _T_1126) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.TinyRocketConfig.fir 208313:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  address = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  d_first_counter = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  opcode_1 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  param_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  size_1 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  source_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sink = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  denied = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inflight = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inflight_opcodes = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  inflight_sizes = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_14[9:0];
  _RAND_15 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_15[9:0];
  _RAND_16 = {1{`RANDOM}};
  watchdog = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_17_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 208519:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 208520:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 208521:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input  [3:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input  [31:0] auto_in_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input  [3:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input  [31:0] auto_in_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output [31:0] auto_in_d_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output [3:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output        auto_out_a_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output [31:0] auto_out_a_bits_address, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output [3:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output [31:0] auto_out_a_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input  [3:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input         auto_out_d_bits_source, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input         auto_out_d_bits_sink, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input  [31:0] auto_out_d_bits_data, // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.TinyRocketConfig.fir 208522:4]
);
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire [3:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [31:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [31:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire  bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [31:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire [31:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire  bundleOut_0_a_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire [1:0] bundleIn_0_d_q_io_enq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire [3:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_enq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_enq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire [31:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_enq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire [3:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_deq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire [31:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
  TLMonitor_45_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.TinyRocketConfig.fir 208529:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_6_inTestHarness bundleOut_0_a_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208556:4]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
  );
  Queue_7_inTestHarness bundleIn_0_d_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.TinyRocketConfig.fir 208570:4]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
    .io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Decoupled.scala 299:17 chipyard.TestHarness.TinyRocketConfig.fir 208568:4]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 208583:4]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 208583:4]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 208569:4]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 208569:4]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 208569:4]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 208569:4]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 208569:4]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 208569:4]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 208569:4]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 208569:4]
  assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 Buffer.scala 37:13 chipyard.TestHarness.TinyRocketConfig.fir 208569:4]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 Decoupled.scala 299:17 chipyard.TestHarness.TinyRocketConfig.fir 208582:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208530:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208531:4]
  assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Decoupled.scala 299:17 chipyard.TestHarness.TinyRocketConfig.fir 208568:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 208583:4]
  assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 208583:4]
  assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 208583:4]
  assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 208583:4]
  assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 208583:4]
  assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 208583:4]
  assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 208583:4]
  assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 Buffer.scala 38:13 chipyard.TestHarness.TinyRocketConfig.fir 208583:4]
  assign bundleOut_0_a_q_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208557:4]
  assign bundleOut_0_a_q_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208558:4]
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 208554:4]
  assign bundleIn_0_d_q_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208571:4]
  assign bundleIn_0_d_q_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208572:4]
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 208554:4]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 208554:4]
  assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 208554:4]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 208554:4]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 208554:4]
  assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 208554:4]
  assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 208554:4]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 208554:4]
  assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.TinyRocketConfig.fir 208552:4 LazyModule.scala 311:12 chipyard.TestHarness.TinyRocketConfig.fir 208554:4]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.TinyRocketConfig.fir 208527:4 LazyModule.scala 309:16 chipyard.TestHarness.TinyRocketConfig.fir 208555:4]
endmodule
module SerialRAM_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 208603:2]
  input         clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 208604:4]
  input         reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 208605:4]
  input         io_ser_in_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  output        io_ser_in_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  output [3:0]  io_ser_in_bits, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  output        io_ser_out_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  input         io_ser_out_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  input  [3:0]  io_ser_out_bits, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  output        io_tsi_ser_in_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  input         io_tsi_ser_in_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  input  [31:0] io_tsi_ser_in_bits, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  input         io_tsi_ser_out_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  output        io_tsi_ser_out_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
  output [31:0] io_tsi_ser_out_bits // @[chipyard.TestHarness.TinyRocketConfig.fir 208607:4]
);
  wire  adapter_clock; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire  adapter_reset; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire  adapter_auto_out_a_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire  adapter_auto_out_a_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire [2:0] adapter_auto_out_a_bits_opcode; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire [3:0] adapter_auto_out_a_bits_size; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire [31:0] adapter_auto_out_a_bits_address; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire [3:0] adapter_auto_out_a_bits_mask; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire [31:0] adapter_auto_out_a_bits_data; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire  adapter_auto_out_d_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire  adapter_auto_out_d_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire [31:0] adapter_auto_out_d_bits_data; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire  adapter_io_serial_in_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire  adapter_io_serial_in_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire [31:0] adapter_io_serial_in_bits; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire  adapter_io_serial_out_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire  adapter_io_serial_out_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire [31:0] adapter_io_serial_out_bits; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
  wire  serdesser_clock; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_reset; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_manager_in_a_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_manager_in_a_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [2:0] serdesser_auto_manager_in_a_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [2:0] serdesser_auto_manager_in_a_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [3:0] serdesser_auto_manager_in_a_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_manager_in_a_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [31:0] serdesser_auto_manager_in_a_bits_address; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [3:0] serdesser_auto_manager_in_a_bits_mask; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [31:0] serdesser_auto_manager_in_a_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_manager_in_a_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_manager_in_d_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_manager_in_d_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [2:0] serdesser_auto_manager_in_d_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [1:0] serdesser_auto_manager_in_d_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [3:0] serdesser_auto_manager_in_d_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_manager_in_d_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_manager_in_d_bits_sink; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_manager_in_d_bits_denied; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [31:0] serdesser_auto_manager_in_d_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_manager_in_d_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_client_out_a_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_client_out_a_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [2:0] serdesser_auto_client_out_a_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [2:0] serdesser_auto_client_out_a_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [2:0] serdesser_auto_client_out_a_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [1:0] serdesser_auto_client_out_a_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [28:0] serdesser_auto_client_out_a_bits_address; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [3:0] serdesser_auto_client_out_a_bits_mask; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [31:0] serdesser_auto_client_out_a_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_client_out_a_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_client_out_d_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_client_out_d_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [2:0] serdesser_auto_client_out_d_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [1:0] serdesser_auto_client_out_d_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [2:0] serdesser_auto_client_out_d_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [1:0] serdesser_auto_client_out_d_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_client_out_d_bits_sink; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_client_out_d_bits_denied; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [31:0] serdesser_auto_client_out_d_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_auto_client_out_d_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_io_ser_in_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_io_ser_in_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [3:0] serdesser_io_ser_in_bits; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_io_ser_out_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  serdesser_io_ser_out_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire [3:0] serdesser_io_ser_out_bits; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
  wire  srams_clock; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire  srams_reset; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire  srams_auto_in_a_ready; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire  srams_auto_in_a_valid; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [2:0] srams_auto_in_a_bits_opcode; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [2:0] srams_auto_in_a_bits_param; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [1:0] srams_auto_in_a_bits_size; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [6:0] srams_auto_in_a_bits_source; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [28:0] srams_auto_in_a_bits_address; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [3:0] srams_auto_in_a_bits_mask; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [31:0] srams_auto_in_a_bits_data; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire  srams_auto_in_a_bits_corrupt; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire  srams_auto_in_d_ready; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire  srams_auto_in_d_valid; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [2:0] srams_auto_in_d_bits_opcode; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [1:0] srams_auto_in_d_bits_size; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [6:0] srams_auto_in_d_bits_source; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire [31:0] srams_auto_in_d_bits_data; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
  wire  xbar_auto_in_a_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_in_a_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [2:0] xbar_auto_in_a_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [2:0] xbar_auto_in_a_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [2:0] xbar_auto_in_a_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [1:0] xbar_auto_in_a_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [28:0] xbar_auto_in_a_bits_address; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [3:0] xbar_auto_in_a_bits_mask; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [31:0] xbar_auto_in_a_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_in_a_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_in_d_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_in_d_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [2:0] xbar_auto_in_d_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [1:0] xbar_auto_in_d_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [2:0] xbar_auto_in_d_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [1:0] xbar_auto_in_d_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_in_d_bits_sink; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_in_d_bits_denied; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [31:0] xbar_auto_in_d_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_in_d_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_out_a_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_out_a_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [2:0] xbar_auto_out_a_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [2:0] xbar_auto_out_a_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [2:0] xbar_auto_out_a_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [1:0] xbar_auto_out_a_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [28:0] xbar_auto_out_a_bits_address; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [3:0] xbar_auto_out_a_bits_mask; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [31:0] xbar_auto_out_a_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_out_a_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_out_d_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_out_d_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [2:0] xbar_auto_out_d_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [1:0] xbar_auto_out_d_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [2:0] xbar_auto_out_d_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [1:0] xbar_auto_out_d_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_out_d_bits_sink; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_out_d_bits_denied; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire [31:0] xbar_auto_out_d_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  xbar_auto_out_d_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
  wire  buffer_clock; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_reset; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [1:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [6:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [28:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [3:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [31:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_in_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [1:0] buffer_auto_in_d_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [1:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [6:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_in_d_bits_sink; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [31:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [1:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [6:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [28:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [3:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [31:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_out_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [1:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [6:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire [31:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [2:0] fragmenter_auto_in_a_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [2:0] fragmenter_auto_in_a_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [1:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [28:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [3:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [31:0] fragmenter_auto_in_a_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_in_a_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [2:0] fragmenter_auto_in_d_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [1:0] fragmenter_auto_in_d_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [1:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_in_d_bits_sink; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_in_d_bits_denied; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [31:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_in_d_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [2:0] fragmenter_auto_out_a_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [2:0] fragmenter_auto_out_a_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [6:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [28:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [3:0] fragmenter_auto_out_a_bits_mask; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [31:0] fragmenter_auto_out_a_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_out_a_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [2:0] fragmenter_auto_out_d_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [1:0] fragmenter_auto_out_d_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [6:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_out_d_bits_sink; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_out_d_bits_denied; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire [31:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  fragmenter_auto_out_d_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
  wire  buffer_1_clock; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_reset; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_in_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_in_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [2:0] buffer_1_auto_in_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [3:0] buffer_1_auto_in_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [31:0] buffer_1_auto_in_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [3:0] buffer_1_auto_in_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [31:0] buffer_1_auto_in_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_in_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_in_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [31:0] buffer_1_auto_in_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_out_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_out_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [2:0] buffer_1_auto_out_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [2:0] buffer_1_auto_out_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [3:0] buffer_1_auto_out_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_out_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [31:0] buffer_1_auto_out_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [3:0] buffer_1_auto_out_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [31:0] buffer_1_auto_out_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_out_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_out_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_out_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [2:0] buffer_1_auto_out_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [1:0] buffer_1_auto_out_d_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [3:0] buffer_1_auto_out_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_out_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_out_d_bits_sink; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_out_d_bits_denied; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire [31:0] buffer_1_auto_out_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  wire  buffer_1_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
  SerialAdapter_inTestHarness adapter ( // @[SerialAdapter.scala 311:27 chipyard.TestHarness.TinyRocketConfig.fir 208613:4]
    .clock(adapter_clock),
    .reset(adapter_reset),
    .auto_out_a_ready(adapter_auto_out_a_ready),
    .auto_out_a_valid(adapter_auto_out_a_valid),
    .auto_out_a_bits_opcode(adapter_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(adapter_auto_out_a_bits_size),
    .auto_out_a_bits_address(adapter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(adapter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(adapter_auto_out_a_bits_data),
    .auto_out_d_ready(adapter_auto_out_d_ready),
    .auto_out_d_valid(adapter_auto_out_d_valid),
    .auto_out_d_bits_data(adapter_auto_out_d_bits_data),
    .io_serial_in_ready(adapter_io_serial_in_ready),
    .io_serial_in_valid(adapter_io_serial_in_valid),
    .io_serial_in_bits(adapter_io_serial_in_bits),
    .io_serial_out_ready(adapter_io_serial_out_ready),
    .io_serial_out_valid(adapter_io_serial_out_valid),
    .io_serial_out_bits(adapter_io_serial_out_bits)
  );
  TLSerdesser_1_inTestHarness serdesser ( // @[SerialAdapter.scala 312:29 chipyard.TestHarness.TinyRocketConfig.fir 208620:4]
    .clock(serdesser_clock),
    .reset(serdesser_reset),
    .auto_manager_in_a_ready(serdesser_auto_manager_in_a_ready),
    .auto_manager_in_a_valid(serdesser_auto_manager_in_a_valid),
    .auto_manager_in_a_bits_opcode(serdesser_auto_manager_in_a_bits_opcode),
    .auto_manager_in_a_bits_param(serdesser_auto_manager_in_a_bits_param),
    .auto_manager_in_a_bits_size(serdesser_auto_manager_in_a_bits_size),
    .auto_manager_in_a_bits_source(serdesser_auto_manager_in_a_bits_source),
    .auto_manager_in_a_bits_address(serdesser_auto_manager_in_a_bits_address),
    .auto_manager_in_a_bits_mask(serdesser_auto_manager_in_a_bits_mask),
    .auto_manager_in_a_bits_data(serdesser_auto_manager_in_a_bits_data),
    .auto_manager_in_a_bits_corrupt(serdesser_auto_manager_in_a_bits_corrupt),
    .auto_manager_in_d_ready(serdesser_auto_manager_in_d_ready),
    .auto_manager_in_d_valid(serdesser_auto_manager_in_d_valid),
    .auto_manager_in_d_bits_opcode(serdesser_auto_manager_in_d_bits_opcode),
    .auto_manager_in_d_bits_param(serdesser_auto_manager_in_d_bits_param),
    .auto_manager_in_d_bits_size(serdesser_auto_manager_in_d_bits_size),
    .auto_manager_in_d_bits_source(serdesser_auto_manager_in_d_bits_source),
    .auto_manager_in_d_bits_sink(serdesser_auto_manager_in_d_bits_sink),
    .auto_manager_in_d_bits_denied(serdesser_auto_manager_in_d_bits_denied),
    .auto_manager_in_d_bits_data(serdesser_auto_manager_in_d_bits_data),
    .auto_manager_in_d_bits_corrupt(serdesser_auto_manager_in_d_bits_corrupt),
    .auto_client_out_a_ready(serdesser_auto_client_out_a_ready),
    .auto_client_out_a_valid(serdesser_auto_client_out_a_valid),
    .auto_client_out_a_bits_opcode(serdesser_auto_client_out_a_bits_opcode),
    .auto_client_out_a_bits_param(serdesser_auto_client_out_a_bits_param),
    .auto_client_out_a_bits_size(serdesser_auto_client_out_a_bits_size),
    .auto_client_out_a_bits_source(serdesser_auto_client_out_a_bits_source),
    .auto_client_out_a_bits_address(serdesser_auto_client_out_a_bits_address),
    .auto_client_out_a_bits_mask(serdesser_auto_client_out_a_bits_mask),
    .auto_client_out_a_bits_data(serdesser_auto_client_out_a_bits_data),
    .auto_client_out_a_bits_corrupt(serdesser_auto_client_out_a_bits_corrupt),
    .auto_client_out_d_ready(serdesser_auto_client_out_d_ready),
    .auto_client_out_d_valid(serdesser_auto_client_out_d_valid),
    .auto_client_out_d_bits_opcode(serdesser_auto_client_out_d_bits_opcode),
    .auto_client_out_d_bits_param(serdesser_auto_client_out_d_bits_param),
    .auto_client_out_d_bits_size(serdesser_auto_client_out_d_bits_size),
    .auto_client_out_d_bits_source(serdesser_auto_client_out_d_bits_source),
    .auto_client_out_d_bits_sink(serdesser_auto_client_out_d_bits_sink),
    .auto_client_out_d_bits_denied(serdesser_auto_client_out_d_bits_denied),
    .auto_client_out_d_bits_data(serdesser_auto_client_out_d_bits_data),
    .auto_client_out_d_bits_corrupt(serdesser_auto_client_out_d_bits_corrupt),
    .io_ser_in_ready(serdesser_io_ser_in_ready),
    .io_ser_in_valid(serdesser_io_ser_in_valid),
    .io_ser_in_bits(serdesser_io_ser_in_bits),
    .io_ser_out_ready(serdesser_io_ser_out_ready),
    .io_ser_out_valid(serdesser_io_ser_out_valid),
    .io_ser_out_bits(serdesser_io_ser_out_bits)
  );
  TLRAM_inTestHarness srams ( // @[SerialAdapter.scala 322:15 chipyard.TestHarness.TinyRocketConfig.fir 208627:4]
    .clock(srams_clock),
    .reset(srams_reset),
    .auto_in_a_ready(srams_auto_in_a_ready),
    .auto_in_a_valid(srams_auto_in_a_valid),
    .auto_in_a_bits_opcode(srams_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(srams_auto_in_a_bits_param),
    .auto_in_a_bits_size(srams_auto_in_a_bits_size),
    .auto_in_a_bits_source(srams_auto_in_a_bits_source),
    .auto_in_a_bits_address(srams_auto_in_a_bits_address),
    .auto_in_a_bits_mask(srams_auto_in_a_bits_mask),
    .auto_in_a_bits_data(srams_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(srams_auto_in_a_bits_corrupt),
    .auto_in_d_ready(srams_auto_in_d_ready),
    .auto_in_d_valid(srams_auto_in_d_valid),
    .auto_in_d_bits_opcode(srams_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(srams_auto_in_d_bits_size),
    .auto_in_d_bits_source(srams_auto_in_d_bits_source),
    .auto_in_d_bits_data(srams_auto_in_d_bits_data)
  );
  TLXbar_9_inTestHarness xbar ( // @[Xbar.scala 142:26 chipyard.TestHarness.TinyRocketConfig.fir 208633:4]
    .auto_in_a_ready(xbar_auto_in_a_ready),
    .auto_in_a_valid(xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(xbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(xbar_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(xbar_auto_in_a_bits_corrupt),
    .auto_in_d_ready(xbar_auto_in_d_ready),
    .auto_in_d_valid(xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(xbar_auto_in_d_bits_param),
    .auto_in_d_bits_size(xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(xbar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(xbar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(xbar_auto_in_d_bits_corrupt),
    .auto_out_a_ready(xbar_auto_out_a_ready),
    .auto_out_a_valid(xbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(xbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(xbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(xbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(xbar_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(xbar_auto_out_a_bits_corrupt),
    .auto_out_d_ready(xbar_auto_out_d_ready),
    .auto_out_d_valid(xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(xbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(xbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(xbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(xbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(xbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(xbar_auto_out_d_bits_corrupt)
  );
  TLBuffer_16_inTestHarness buffer ( // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208639:4]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data)
  );
  TLFragmenter_8_inTestHarness fragmenter ( // @[Fragmenter.scala 333:34 chipyard.TestHarness.TinyRocketConfig.fir 208645:4]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(fragmenter_auto_in_d_bits_param),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_sink(fragmenter_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(fragmenter_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fragmenter_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(fragmenter_auto_out_d_bits_param),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_sink(fragmenter_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(fragmenter_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fragmenter_auto_out_d_bits_corrupt)
  );
  TLBuffer_17_inTestHarness buffer_1 ( // @[Buffer.scala 68:28 chipyard.TestHarness.TinyRocketConfig.fir 208651:4]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_a_ready(buffer_1_auto_in_a_ready),
    .auto_in_a_valid(buffer_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
    .auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_1_auto_in_d_ready),
    .auto_in_d_valid(buffer_1_auto_in_d_valid),
    .auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
    .auto_out_a_ready(buffer_1_auto_out_a_ready),
    .auto_out_a_valid(buffer_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_1_auto_out_a_bits_corrupt),
    .auto_out_d_ready(buffer_1_auto_out_d_ready),
    .auto_out_d_valid(buffer_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
  );
  assign io_ser_in_valid = serdesser_io_ser_out_valid; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.TinyRocketConfig.fir 208667:4]
  assign io_ser_in_bits = serdesser_io_ser_out_bits; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.TinyRocketConfig.fir 208666:4]
  assign io_ser_out_ready = serdesser_io_ser_in_ready; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.TinyRocketConfig.fir 208665:4]
  assign io_tsi_ser_in_ready = adapter_io_serial_in_ready; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.TinyRocketConfig.fir 208674:4]
  assign io_tsi_ser_out_valid = adapter_io_serial_out_valid; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.TinyRocketConfig.fir 208670:4]
  assign io_tsi_ser_out_bits = adapter_io_serial_out_bits; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.TinyRocketConfig.fir 208669:4]
  assign adapter_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208618:4]
  assign adapter_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208619:4]
  assign adapter_auto_out_a_ready = buffer_1_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208657:4]
  assign adapter_auto_out_d_valid = buffer_1_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208657:4]
  assign adapter_auto_out_d_bits_data = buffer_1_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208657:4]
  assign adapter_io_serial_in_valid = io_tsi_ser_in_valid; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.TinyRocketConfig.fir 208673:4]
  assign adapter_io_serial_in_bits = io_tsi_ser_in_bits; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.TinyRocketConfig.fir 208672:4]
  assign adapter_io_serial_out_ready = io_tsi_ser_out_ready; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.TinyRocketConfig.fir 208671:4]
  assign serdesser_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208625:4]
  assign serdesser_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208626:4]
  assign serdesser_auto_manager_in_a_valid = buffer_1_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign serdesser_auto_manager_in_a_bits_opcode = buffer_1_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign serdesser_auto_manager_in_a_bits_param = buffer_1_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign serdesser_auto_manager_in_a_bits_size = buffer_1_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign serdesser_auto_manager_in_a_bits_source = buffer_1_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign serdesser_auto_manager_in_a_bits_address = buffer_1_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign serdesser_auto_manager_in_a_bits_mask = buffer_1_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign serdesser_auto_manager_in_a_bits_data = buffer_1_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign serdesser_auto_manager_in_a_bits_corrupt = buffer_1_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign serdesser_auto_manager_in_d_ready = buffer_1_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign serdesser_auto_client_out_a_ready = xbar_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign serdesser_auto_client_out_d_valid = xbar_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign serdesser_auto_client_out_d_bits_opcode = xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign serdesser_auto_client_out_d_bits_param = xbar_auto_in_d_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign serdesser_auto_client_out_d_bits_size = xbar_auto_in_d_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign serdesser_auto_client_out_d_bits_source = xbar_auto_in_d_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign serdesser_auto_client_out_d_bits_sink = xbar_auto_in_d_bits_sink; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign serdesser_auto_client_out_d_bits_denied = xbar_auto_in_d_bits_denied; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign serdesser_auto_client_out_d_bits_data = xbar_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign serdesser_auto_client_out_d_bits_corrupt = xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign serdesser_io_ser_in_valid = io_ser_out_valid; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.TinyRocketConfig.fir 208664:4]
  assign serdesser_io_ser_in_bits = io_ser_out_bits; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.TinyRocketConfig.fir 208663:4]
  assign serdesser_io_ser_out_ready = io_ser_in_ready; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.TinyRocketConfig.fir 208668:4]
  assign srams_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208631:4]
  assign srams_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208632:4]
  assign srams_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign srams_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign srams_auto_in_a_bits_param = buffer_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign srams_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign srams_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign srams_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign srams_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign srams_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign srams_auto_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign srams_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign xbar_auto_in_a_valid = serdesser_auto_client_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign xbar_auto_in_a_bits_opcode = serdesser_auto_client_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign xbar_auto_in_a_bits_param = serdesser_auto_client_out_a_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign xbar_auto_in_a_bits_size = serdesser_auto_client_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign xbar_auto_in_a_bits_source = serdesser_auto_client_out_a_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign xbar_auto_in_a_bits_address = serdesser_auto_client_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign xbar_auto_in_a_bits_mask = serdesser_auto_client_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign xbar_auto_in_a_bits_data = serdesser_auto_client_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign xbar_auto_in_a_bits_corrupt = serdesser_auto_client_out_a_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign xbar_auto_in_d_ready = serdesser_auto_client_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208658:4]
  assign xbar_auto_out_a_ready = fragmenter_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign xbar_auto_out_d_valid = fragmenter_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign xbar_auto_out_d_bits_opcode = fragmenter_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign xbar_auto_out_d_bits_param = fragmenter_auto_in_d_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign xbar_auto_out_d_bits_size = fragmenter_auto_in_d_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign xbar_auto_out_d_bits_source = fragmenter_auto_in_d_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign xbar_auto_out_d_bits_sink = fragmenter_auto_in_d_bits_sink; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign xbar_auto_out_d_bits_denied = fragmenter_auto_in_d_bits_denied; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign xbar_auto_out_d_bits_data = fragmenter_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign xbar_auto_out_d_bits_corrupt = fragmenter_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign buffer_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208643:4]
  assign buffer_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208644:4]
  assign buffer_auto_in_a_valid = fragmenter_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_auto_in_a_bits_opcode = fragmenter_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_auto_in_a_bits_param = fragmenter_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_auto_in_a_bits_size = fragmenter_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_auto_in_a_bits_source = fragmenter_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_auto_in_a_bits_address = fragmenter_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_auto_in_a_bits_mask = fragmenter_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_auto_in_a_bits_data = fragmenter_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_auto_in_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_auto_in_d_ready = fragmenter_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_auto_out_a_ready = srams_auto_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign buffer_auto_out_d_valid = srams_auto_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign buffer_auto_out_d_bits_opcode = srams_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign buffer_auto_out_d_bits_size = srams_auto_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign buffer_auto_out_d_bits_source = srams_auto_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign buffer_auto_out_d_bits_data = srams_auto_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208660:4]
  assign fragmenter_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208649:4]
  assign fragmenter_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208650:4]
  assign fragmenter_auto_in_a_valid = xbar_auto_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign fragmenter_auto_in_a_bits_opcode = xbar_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign fragmenter_auto_in_a_bits_param = xbar_auto_out_a_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign fragmenter_auto_in_a_bits_size = xbar_auto_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign fragmenter_auto_in_a_bits_source = xbar_auto_out_a_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign fragmenter_auto_in_a_bits_address = xbar_auto_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign fragmenter_auto_in_a_bits_mask = xbar_auto_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign fragmenter_auto_in_a_bits_data = xbar_auto_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign fragmenter_auto_in_a_bits_corrupt = xbar_auto_out_a_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign fragmenter_auto_in_d_ready = xbar_auto_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208659:4]
  assign fragmenter_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign fragmenter_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign fragmenter_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign fragmenter_auto_out_d_bits_param = buffer_auto_in_d_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign fragmenter_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign fragmenter_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign fragmenter_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign fragmenter_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign fragmenter_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign fragmenter_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208661:4]
  assign buffer_1_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208655:4]
  assign buffer_1_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208656:4]
  assign buffer_1_auto_in_a_valid = adapter_auto_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208657:4]
  assign buffer_1_auto_in_a_bits_opcode = adapter_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208657:4]
  assign buffer_1_auto_in_a_bits_size = adapter_auto_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208657:4]
  assign buffer_1_auto_in_a_bits_address = adapter_auto_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208657:4]
  assign buffer_1_auto_in_a_bits_mask = adapter_auto_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208657:4]
  assign buffer_1_auto_in_a_bits_data = adapter_auto_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208657:4]
  assign buffer_1_auto_in_d_ready = adapter_auto_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.TinyRocketConfig.fir 208657:4]
  assign buffer_1_auto_out_a_ready = serdesser_auto_manager_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign buffer_1_auto_out_d_valid = serdesser_auto_manager_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign buffer_1_auto_out_d_bits_opcode = serdesser_auto_manager_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign buffer_1_auto_out_d_bits_param = serdesser_auto_manager_in_d_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign buffer_1_auto_out_d_bits_size = serdesser_auto_manager_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign buffer_1_auto_out_d_bits_source = serdesser_auto_manager_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign buffer_1_auto_out_d_bits_sink = serdesser_auto_manager_in_d_bits_sink; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign buffer_1_auto_out_d_bits_denied = serdesser_auto_manager_in_d_bits_denied; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign buffer_1_auto_out_d_bits_data = serdesser_auto_manager_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
  assign buffer_1_auto_out_d_bits_corrupt = serdesser_auto_manager_in_d_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.TinyRocketConfig.fir 208662:4]
endmodule
module Queue_26_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 208685:2]
  input        clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 208686:4]
  input        reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 208687:4]
  output       io_enq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 208688:4]
  input        io_enq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 208688:4]
  input  [7:0] io_enq_bits, // @[chipyard.TestHarness.TinyRocketConfig.fir 208688:4]
  input        io_deq_ready, // @[chipyard.TestHarness.TinyRocketConfig.fir 208688:4]
  output       io_deq_valid, // @[chipyard.TestHarness.TinyRocketConfig.fir 208688:4]
  output [7:0] io_deq_bits // @[chipyard.TestHarness.TinyRocketConfig.fir 208688:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:127]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 208690:4]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 208690:4]
  wire [6:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 208690:4]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 208690:4]
  wire [6:0] ram_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 208690:4]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 208690:4]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 208690:4]
  reg [6:0] enq_ptr_value; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208691:4]
  reg [6:0] deq_ptr_value; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208692:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 208693:4]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33 chipyard.TestHarness.TinyRocketConfig.fir 208694:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.TinyRocketConfig.fir 208695:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.TinyRocketConfig.fir 208696:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.TinyRocketConfig.fir 208697:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 208698:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.TinyRocketConfig.fir 208701:4]
  wire [6:0] _value_T_1 = enq_ptr_value + 7'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 208709:6]
  wire [6:0] _value_T_3 = deq_ptr_value + 7'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 208715:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.TinyRocketConfig.fir 208718:4]
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 208690:4]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.TinyRocketConfig.fir 208724:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.TinyRocketConfig.fir 208722:4]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.TinyRocketConfig.fir 208727:4]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.TinyRocketConfig.fir 208690:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208691:4]
      enq_ptr_value <= 7'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208691:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.TinyRocketConfig.fir 208704:4]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 208710:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208692:4]
      deq_ptr_value <= 7'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208692:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.TinyRocketConfig.fir 208712:4]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 208716:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 208693:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.TinyRocketConfig.fir 208693:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.TinyRocketConfig.fir 208719:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.TinyRocketConfig.fir 208720:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module UARTAdapter_inTestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 208793:2]
  input   clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 208794:4]
  input   reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 208795:4]
  input   io_uart_txd, // @[chipyard.TestHarness.TinyRocketConfig.fir 208796:4]
  output  io_uart_rxd // @[chipyard.TestHarness.TinyRocketConfig.fir 208796:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  txfifo_clock; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.TinyRocketConfig.fir 208798:4]
  wire  txfifo_reset; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.TinyRocketConfig.fir 208798:4]
  wire  txfifo_io_enq_ready; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.TinyRocketConfig.fir 208798:4]
  wire  txfifo_io_enq_valid; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.TinyRocketConfig.fir 208798:4]
  wire [7:0] txfifo_io_enq_bits; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.TinyRocketConfig.fir 208798:4]
  wire  txfifo_io_deq_ready; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.TinyRocketConfig.fir 208798:4]
  wire  txfifo_io_deq_valid; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.TinyRocketConfig.fir 208798:4]
  wire [7:0] txfifo_io_deq_bits; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.TinyRocketConfig.fir 208798:4]
  wire  rxfifo_clock; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.TinyRocketConfig.fir 208801:4]
  wire  rxfifo_reset; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.TinyRocketConfig.fir 208801:4]
  wire  rxfifo_io_enq_ready; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.TinyRocketConfig.fir 208801:4]
  wire  rxfifo_io_enq_valid; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.TinyRocketConfig.fir 208801:4]
  wire [7:0] rxfifo_io_enq_bits; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.TinyRocketConfig.fir 208801:4]
  wire  rxfifo_io_deq_ready; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.TinyRocketConfig.fir 208801:4]
  wire  rxfifo_io_deq_valid; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.TinyRocketConfig.fir 208801:4]
  wire [7:0] rxfifo_io_deq_bits; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.TinyRocketConfig.fir 208801:4]
  wire  sim_clock; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.TinyRocketConfig.fir 208950:4]
  wire  sim_reset; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.TinyRocketConfig.fir 208950:4]
  wire  sim_serial_in_ready; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.TinyRocketConfig.fir 208950:4]
  wire  sim_serial_in_valid; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.TinyRocketConfig.fir 208950:4]
  wire [7:0] sim_serial_in_bits; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.TinyRocketConfig.fir 208950:4]
  wire  sim_serial_out_ready; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.TinyRocketConfig.fir 208950:4]
  wire  sim_serial_out_valid; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.TinyRocketConfig.fir 208950:4]
  wire [7:0] sim_serial_out_bits; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.TinyRocketConfig.fir 208950:4]
  reg [1:0] txState; // @[UARTAdapter.scala 38:24 chipyard.TestHarness.TinyRocketConfig.fir 208804:4]
  reg [7:0] txData; // @[UARTAdapter.scala 39:19 chipyard.TestHarness.TinyRocketConfig.fir 208805:4]
  wire  _T = txState == 2'h2; // @[UARTAdapter.scala 41:49 chipyard.TestHarness.TinyRocketConfig.fir 208806:4]
  wire  _T_1 = _T & txfifo_io_enq_ready; // @[UARTAdapter.scala 41:61 chipyard.TestHarness.TinyRocketConfig.fir 208807:4]
  reg [2:0] txDataIdx; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208808:4]
  wire  wrap_wrap = txDataIdx == 3'h7; // @[Counter.scala 72:24 chipyard.TestHarness.TinyRocketConfig.fir 208812:6]
  wire [2:0] _wrap_value_T_1 = txDataIdx + 3'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 208814:6]
  wire  txDataWrap = _T_1 & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208811:4 Counter.scala 118:24 chipyard.TestHarness.TinyRocketConfig.fir 208816:6 chipyard.TestHarness.TinyRocketConfig.fir 208810:4]
  wire  _T_2 = txState == 2'h1; // @[UARTAdapter.scala 43:51 chipyard.TestHarness.TinyRocketConfig.fir 208818:4]
  wire  _T_3 = _T_2 & txfifo_io_enq_ready; // @[UARTAdapter.scala 43:63 chipyard.TestHarness.TinyRocketConfig.fir 208819:4]
  reg [9:0] txBaudCount; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208820:4]
  wire  wrap_wrap_1 = txBaudCount == 10'h363; // @[Counter.scala 72:24 chipyard.TestHarness.TinyRocketConfig.fir 208824:6]
  wire [9:0] _wrap_value_T_3 = txBaudCount + 10'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 208826:6]
  wire  txBaudWrap = _T_3 & wrap_wrap_1; // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208823:4 Counter.scala 118:24 chipyard.TestHarness.TinyRocketConfig.fir 208831:6 chipyard.TestHarness.TinyRocketConfig.fir 208822:4]
  wire  _T_4 = txState == 2'h0; // @[UARTAdapter.scala 44:53 chipyard.TestHarness.TinyRocketConfig.fir 208833:4]
  wire  _T_5 = ~io_uart_txd; // @[UARTAdapter.scala 44:80 chipyard.TestHarness.TinyRocketConfig.fir 208834:4]
  wire  _T_6 = _T_4 & _T_5; // @[UARTAdapter.scala 44:65 chipyard.TestHarness.TinyRocketConfig.fir 208835:4]
  wire  _T_7 = _T_6 & txfifo_io_enq_ready; // @[UARTAdapter.scala 44:88 chipyard.TestHarness.TinyRocketConfig.fir 208836:4]
  reg [1:0] txSlackCount; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208837:4]
  wire  wrap_wrap_2 = txSlackCount == 2'h3; // @[Counter.scala 72:24 chipyard.TestHarness.TinyRocketConfig.fir 208841:6]
  wire [1:0] _wrap_value_T_5 = txSlackCount + 2'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 208843:6]
  wire  txSlackWrap = _T_7 & wrap_wrap_2; // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208840:4 Counter.scala 118:24 chipyard.TestHarness.TinyRocketConfig.fir 208845:6 chipyard.TestHarness.TinyRocketConfig.fir 208839:4]
  wire  _T_8 = 2'h0 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.TinyRocketConfig.fir 208847:4]
  wire  _T_9 = 2'h1 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.TinyRocketConfig.fir 208855:6]
  wire  _T_10 = 2'h2 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.TinyRocketConfig.fir 208862:8]
  wire [7:0] _GEN_35 = {{7'd0}, io_uart_txd}; // @[UARTAdapter.scala 60:41 chipyard.TestHarness.TinyRocketConfig.fir 208865:12]
  wire [7:0] _txData_T = _GEN_35 << txDataIdx; // @[UARTAdapter.scala 60:41 chipyard.TestHarness.TinyRocketConfig.fir 208865:12]
  wire [7:0] _txData_T_1 = txData | _txData_T; // @[UARTAdapter.scala 60:26 chipyard.TestHarness.TinyRocketConfig.fir 208866:12]
  wire [1:0] _txState_T_1 = io_uart_txd ? 2'h0 : 2'h3; // @[UARTAdapter.scala 63:23 chipyard.TestHarness.TinyRocketConfig.fir 208871:12]
  wire [1:0] _GEN_11 = txfifo_io_enq_ready ? 2'h1 : txState; // @[UARTAdapter.scala 64:39 chipyard.TestHarness.TinyRocketConfig.fir 208875:12 UARTAdapter.scala 65:17 chipyard.TestHarness.TinyRocketConfig.fir 208876:14 UARTAdapter.scala 38:24 chipyard.TestHarness.TinyRocketConfig.fir 208804:4]
  wire [1:0] _GEN_12 = txDataWrap ? _txState_T_1 : _GEN_11; // @[UARTAdapter.scala 62:24 chipyard.TestHarness.TinyRocketConfig.fir 208869:10 UARTAdapter.scala 63:17 chipyard.TestHarness.TinyRocketConfig.fir 208872:12]
  wire  _T_11 = 2'h3 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.TinyRocketConfig.fir 208880:10]
  wire  _T_13 = io_uart_txd & txfifo_io_enq_ready; // @[UARTAdapter.scala 69:32 chipyard.TestHarness.TinyRocketConfig.fir 208883:12]
  wire [1:0] _GEN_13 = _T_13 ? 2'h0 : txState; // @[UARTAdapter.scala 69:56 chipyard.TestHarness.TinyRocketConfig.fir 208884:12 UARTAdapter.scala 70:17 chipyard.TestHarness.TinyRocketConfig.fir 208885:14 UARTAdapter.scala 38:24 chipyard.TestHarness.TinyRocketConfig.fir 208804:4]
  wire [1:0] _GEN_14 = _T_11 ? _GEN_13 : txState; // @[Conditional.scala 39:67 chipyard.TestHarness.TinyRocketConfig.fir 208881:10 UARTAdapter.scala 38:24 chipyard.TestHarness.TinyRocketConfig.fir 208804:4]
  reg [1:0] rxState; // @[UARTAdapter.scala 79:24 chipyard.TestHarness.TinyRocketConfig.fir 208890:4]
  reg [9:0] rxBaudCount; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208891:4]
  wire  wrap_wrap_3 = rxBaudCount == 10'h363; // @[Counter.scala 72:24 chipyard.TestHarness.TinyRocketConfig.fir 208895:6]
  wire [9:0] _wrap_value_T_7 = rxBaudCount + 10'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 208897:6]
  wire  rxBaudWrap = txfifo_io_enq_ready & wrap_wrap_3; // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208894:4 Counter.scala 118:24 chipyard.TestHarness.TinyRocketConfig.fir 208902:6 chipyard.TestHarness.TinyRocketConfig.fir 208893:4]
  wire  _T_14 = rxState == 2'h2; // @[UARTAdapter.scala 83:49 chipyard.TestHarness.TinyRocketConfig.fir 208904:4]
  wire  _T_15 = _T_14 & txfifo_io_enq_ready; // @[UARTAdapter.scala 83:61 chipyard.TestHarness.TinyRocketConfig.fir 208905:4]
  wire  _T_16 = _T_15 & rxBaudWrap; // @[UARTAdapter.scala 83:84 chipyard.TestHarness.TinyRocketConfig.fir 208906:4]
  reg [2:0] rxDataIdx; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208907:4]
  wire  wrap_wrap_4 = rxDataIdx == 3'h7; // @[Counter.scala 72:24 chipyard.TestHarness.TinyRocketConfig.fir 208911:6]
  wire [2:0] _wrap_value_T_9 = rxDataIdx + 3'h1; // @[Counter.scala 76:24 chipyard.TestHarness.TinyRocketConfig.fir 208913:6]
  wire  rxDataWrap = _T_16 & wrap_wrap_4; // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208910:4 Counter.scala 118:24 chipyard.TestHarness.TinyRocketConfig.fir 208915:6 chipyard.TestHarness.TinyRocketConfig.fir 208909:4]
  wire  _T_17 = 2'h0 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.TinyRocketConfig.fir 208918:4]
  wire  _T_18 = rxBaudWrap & rxfifo_io_deq_valid; // @[UARTAdapter.scala 89:24 chipyard.TestHarness.TinyRocketConfig.fir 208921:6]
  wire  _T_19 = 2'h1 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.TinyRocketConfig.fir 208927:6]
  wire  _T_20 = 2'h2 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.TinyRocketConfig.fir 208935:8]
  wire [7:0] _io_uart_rxd_T = rxfifo_io_deq_bits >> rxDataIdx; // @[UARTAdapter.scala 100:42 chipyard.TestHarness.TinyRocketConfig.fir 208937:10]
  wire  _T_21 = rxDataWrap & rxBaudWrap; // @[UARTAdapter.scala 101:23 chipyard.TestHarness.TinyRocketConfig.fir 208940:10]
  wire [1:0] _GEN_28 = _T_21 ? 2'h0 : rxState; // @[UARTAdapter.scala 101:38 chipyard.TestHarness.TinyRocketConfig.fir 208941:10 UARTAdapter.scala 102:17 chipyard.TestHarness.TinyRocketConfig.fir 208942:12 UARTAdapter.scala 79:24 chipyard.TestHarness.TinyRocketConfig.fir 208890:4]
  wire  _GEN_29 = _T_20 ? _io_uart_rxd_T[0] : 1'h1; // @[Conditional.scala 39:67 chipyard.TestHarness.TinyRocketConfig.fir 208936:8 UARTAdapter.scala 100:19 chipyard.TestHarness.TinyRocketConfig.fir 208939:10 UARTAdapter.scala 85:15 chipyard.TestHarness.TinyRocketConfig.fir 208917:4]
  wire  _GEN_31 = _T_19 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67 chipyard.TestHarness.TinyRocketConfig.fir 208928:6 UARTAdapter.scala 94:19 chipyard.TestHarness.TinyRocketConfig.fir 208929:8]
  wire  _rxfifo_io_deq_ready_T_1 = _T_14 & rxDataWrap; // @[UARTAdapter.scala 106:48 chipyard.TestHarness.TinyRocketConfig.fir 208946:4]
  wire  _rxfifo_io_deq_ready_T_2 = _rxfifo_io_deq_ready_T_1 & rxBaudWrap; // @[UARTAdapter.scala 106:62 chipyard.TestHarness.TinyRocketConfig.fir 208947:4]
  Queue_26_inTestHarness txfifo ( // @[UARTAdapter.scala 32:22 chipyard.TestHarness.TinyRocketConfig.fir 208798:4]
    .clock(txfifo_clock),
    .reset(txfifo_reset),
    .io_enq_ready(txfifo_io_enq_ready),
    .io_enq_valid(txfifo_io_enq_valid),
    .io_enq_bits(txfifo_io_enq_bits),
    .io_deq_ready(txfifo_io_deq_ready),
    .io_deq_valid(txfifo_io_deq_valid),
    .io_deq_bits(txfifo_io_deq_bits)
  );
  Queue_26_inTestHarness rxfifo ( // @[UARTAdapter.scala 33:22 chipyard.TestHarness.TinyRocketConfig.fir 208801:4]
    .clock(rxfifo_clock),
    .reset(rxfifo_reset),
    .io_enq_ready(rxfifo_io_enq_ready),
    .io_enq_valid(rxfifo_io_enq_valid),
    .io_enq_bits(rxfifo_io_enq_bits),
    .io_deq_ready(rxfifo_io_deq_ready),
    .io_deq_valid(rxfifo_io_deq_valid),
    .io_deq_bits(rxfifo_io_deq_bits)
  );
  SimUART #(.UARTNO(0)) sim ( // @[UARTAdapter.scala 108:19 chipyard.TestHarness.TinyRocketConfig.fir 208950:4]
    .clock(sim_clock),
    .reset(sim_reset),
    .serial_in_ready(sim_serial_in_ready),
    .serial_in_valid(sim_serial_in_valid),
    .serial_in_bits(sim_serial_in_bits),
    .serial_out_ready(sim_serial_out_ready),
    .serial_out_valid(sim_serial_out_valid),
    .serial_out_bits(sim_serial_out_bits)
  );
  assign io_uart_rxd = _T_17 | _GEN_31; // @[Conditional.scala 40:58 chipyard.TestHarness.TinyRocketConfig.fir 208919:4 UARTAdapter.scala 88:19 chipyard.TestHarness.TinyRocketConfig.fir 208920:6]
  assign txfifo_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208799:4]
  assign txfifo_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208800:4]
  assign txfifo_io_enq_valid = _T_1 & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208811:4 Counter.scala 118:24 chipyard.TestHarness.TinyRocketConfig.fir 208816:6 chipyard.TestHarness.TinyRocketConfig.fir 208810:4]
  assign txfifo_io_enq_bits = txData; // @[UARTAdapter.scala 75:23 chipyard.TestHarness.TinyRocketConfig.fir 208888:4]
  assign txfifo_io_deq_ready = sim_serial_out_ready; // @[UARTAdapter.scala 115:23 chipyard.TestHarness.TinyRocketConfig.fir 208959:4]
  assign rxfifo_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 208802:4]
  assign rxfifo_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208803:4]
  assign rxfifo_io_enq_valid = sim_serial_in_valid; // @[UARTAdapter.scala 118:23 chipyard.TestHarness.TinyRocketConfig.fir 208961:4]
  assign rxfifo_io_enq_bits = sim_serial_in_bits; // @[UARTAdapter.scala 117:22 chipyard.TestHarness.TinyRocketConfig.fir 208960:4]
  assign rxfifo_io_deq_ready = _rxfifo_io_deq_ready_T_2 & txfifo_io_enq_ready; // @[UARTAdapter.scala 106:76 chipyard.TestHarness.TinyRocketConfig.fir 208948:4]
  assign sim_clock = clock; // @[UARTAdapter.scala 110:16 chipyard.TestHarness.TinyRocketConfig.fir 208954:4]
  assign sim_reset = reset; // @[UARTAdapter.scala 111:25 chipyard.TestHarness.TinyRocketConfig.fir 208955:4]
  assign sim_serial_in_ready = rxfifo_io_enq_ready; // @[UARTAdapter.scala 119:26 chipyard.TestHarness.TinyRocketConfig.fir 208962:4]
  assign sim_serial_out_valid = txfifo_io_deq_valid; // @[UARTAdapter.scala 114:27 chipyard.TestHarness.TinyRocketConfig.fir 208958:4]
  assign sim_serial_out_bits = txfifo_io_deq_bits; // @[UARTAdapter.scala 113:26 chipyard.TestHarness.TinyRocketConfig.fir 208957:4]
  always @(posedge clock) begin
    if (reset) begin // @[UARTAdapter.scala 38:24 chipyard.TestHarness.TinyRocketConfig.fir 208804:4]
      txState <= 2'h0; // @[UARTAdapter.scala 38:24 chipyard.TestHarness.TinyRocketConfig.fir 208804:4]
    end else if (_T_8) begin // @[Conditional.scala 40:58 chipyard.TestHarness.TinyRocketConfig.fir 208848:4]
      if (txSlackWrap) begin // @[UARTAdapter.scala 48:25 chipyard.TestHarness.TinyRocketConfig.fir 208849:6]
        txState <= 2'h1; // @[UARTAdapter.scala 50:17 chipyard.TestHarness.TinyRocketConfig.fir 208851:8]
      end
    end else if (_T_9) begin // @[Conditional.scala 39:67 chipyard.TestHarness.TinyRocketConfig.fir 208856:6]
      if (txBaudWrap) begin // @[UARTAdapter.scala 54:24 chipyard.TestHarness.TinyRocketConfig.fir 208857:8]
        txState <= 2'h2; // @[UARTAdapter.scala 55:17 chipyard.TestHarness.TinyRocketConfig.fir 208858:10]
      end
    end else if (_T_10) begin // @[Conditional.scala 39:67 chipyard.TestHarness.TinyRocketConfig.fir 208863:8]
      txState <= _GEN_12;
    end else begin
      txState <= _GEN_14;
    end
    if (_T_8) begin // @[Conditional.scala 40:58 chipyard.TestHarness.TinyRocketConfig.fir 208848:4]
      if (txSlackWrap) begin // @[UARTAdapter.scala 48:25 chipyard.TestHarness.TinyRocketConfig.fir 208849:6]
        txData <= 8'h0; // @[UARTAdapter.scala 49:17 chipyard.TestHarness.TinyRocketConfig.fir 208850:8]
      end
    end else if (!(_T_9)) begin // @[Conditional.scala 39:67 chipyard.TestHarness.TinyRocketConfig.fir 208856:6]
      if (_T_10) begin // @[Conditional.scala 39:67 chipyard.TestHarness.TinyRocketConfig.fir 208863:8]
        if (txfifo_io_enq_ready) begin // @[UARTAdapter.scala 59:34 chipyard.TestHarness.TinyRocketConfig.fir 208864:10]
          txData <= _txData_T_1; // @[UARTAdapter.scala 60:16 chipyard.TestHarness.TinyRocketConfig.fir 208867:12]
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208808:4]
      txDataIdx <= 3'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208808:4]
    end else if (_T_1) begin // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208811:4]
      txDataIdx <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 208815:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208820:4]
      txBaudCount <= 10'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208820:4]
    end else if (_T_3) begin // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208823:4]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20 chipyard.TestHarness.TinyRocketConfig.fir 208828:6]
        txBaudCount <= 10'h0; // @[Counter.scala 86:28 chipyard.TestHarness.TinyRocketConfig.fir 208829:8]
      end else begin
        txBaudCount <= _wrap_value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 208827:6]
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208837:4]
      txSlackCount <= 2'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208837:4]
    end else if (_T_7) begin // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208840:4]
      txSlackCount <= _wrap_value_T_5; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 208844:6]
    end
    if (reset) begin // @[UARTAdapter.scala 79:24 chipyard.TestHarness.TinyRocketConfig.fir 208890:4]
      rxState <= 2'h0; // @[UARTAdapter.scala 79:24 chipyard.TestHarness.TinyRocketConfig.fir 208890:4]
    end else if (_T_17) begin // @[Conditional.scala 40:58 chipyard.TestHarness.TinyRocketConfig.fir 208919:4]
      if (_T_18) begin // @[UARTAdapter.scala 89:48 chipyard.TestHarness.TinyRocketConfig.fir 208922:6]
        rxState <= 2'h1; // @[UARTAdapter.scala 90:17 chipyard.TestHarness.TinyRocketConfig.fir 208923:8]
      end
    end else if (_T_19) begin // @[Conditional.scala 39:67 chipyard.TestHarness.TinyRocketConfig.fir 208928:6]
      if (rxBaudWrap) begin // @[UARTAdapter.scala 95:24 chipyard.TestHarness.TinyRocketConfig.fir 208930:8]
        rxState <= 2'h2; // @[UARTAdapter.scala 96:17 chipyard.TestHarness.TinyRocketConfig.fir 208931:10]
      end
    end else if (_T_20) begin // @[Conditional.scala 39:67 chipyard.TestHarness.TinyRocketConfig.fir 208936:8]
      rxState <= _GEN_28;
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208891:4]
      rxBaudCount <= 10'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208891:4]
    end else if (txfifo_io_enq_ready) begin // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208894:4]
      if (wrap_wrap_3) begin // @[Counter.scala 86:20 chipyard.TestHarness.TinyRocketConfig.fir 208899:6]
        rxBaudCount <= 10'h0; // @[Counter.scala 86:28 chipyard.TestHarness.TinyRocketConfig.fir 208900:8]
      end else begin
        rxBaudCount <= _wrap_value_T_7; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 208898:6]
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208907:4]
      rxDataIdx <= 3'h0; // @[Counter.scala 60:40 chipyard.TestHarness.TinyRocketConfig.fir 208907:4]
    end else if (_T_16) begin // @[Counter.scala 118:17 chipyard.TestHarness.TinyRocketConfig.fir 208910:4]
      rxDataIdx <= _wrap_value_T_9; // @[Counter.scala 76:15 chipyard.TestHarness.TinyRocketConfig.fir 208914:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  txState = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  txData = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  txDataIdx = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  txBaudCount = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  txSlackCount = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  rxState = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  rxBaudCount = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  rxDataIdx = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TestHarness( // @[chipyard.TestHarness.TinyRocketConfig.fir 208964:2]
  input   clock, // @[chipyard.TestHarness.TinyRocketConfig.fir 208965:4]
  input   reset, // @[chipyard.TestHarness.TinyRocketConfig.fir 208966:4]
  output  io_success // @[chipyard.TestHarness.TinyRocketConfig.fir 208967:4]
);
  wire  chiptop_jtag_TCK; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_jtag_TMS; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_jtag_TDI; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_jtag_TDO_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_jtag_TDO_driven; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_serial_tl_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_serial_tl_bits_in_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_serial_tl_bits_in_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire [3:0] chiptop_serial_tl_bits_in_bits; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_serial_tl_bits_out_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_serial_tl_bits_out_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire [3:0] chiptop_serial_tl_bits_out_bits; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_uart_0_txd; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_uart_0_rxd; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_reset_wire_reset; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  chiptop_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
  wire  SimJTAG_clock; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire  SimJTAG_reset; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire  SimJTAG_jtag_TRSTn; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire  SimJTAG_jtag_TCK; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire  SimJTAG_jtag_TMS; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire  SimJTAG_jtag_TDI; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire  SimJTAG_jtag_TDO_data; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire  SimJTAG_jtag_TDO_driven; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire  SimJTAG_enable; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire  SimJTAG_init_done; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire [31:0] SimJTAG_exit; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 208998:4]
  wire  ram_clock; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire  ram_reset; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire  ram_io_ser_in_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire  ram_io_ser_in_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire [3:0] ram_io_ser_in_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire  ram_io_ser_out_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire  ram_io_ser_out_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire [3:0] ram_io_ser_out_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire  ram_io_tsi_ser_in_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire  ram_io_tsi_ser_in_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire [31:0] ram_io_tsi_ser_in_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire  ram_io_tsi_ser_out_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire  ram_io_tsi_ser_out_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire [31:0] ram_io_tsi_ser_out_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
  wire  success_sim_clock; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.TinyRocketConfig.fir 209028:4]
  wire  success_sim_reset; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.TinyRocketConfig.fir 209028:4]
  wire  success_sim_serial_in_ready; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.TinyRocketConfig.fir 209028:4]
  wire  success_sim_serial_in_valid; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.TinyRocketConfig.fir 209028:4]
  wire [31:0] success_sim_serial_in_bits; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.TinyRocketConfig.fir 209028:4]
  wire  success_sim_serial_out_ready; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.TinyRocketConfig.fir 209028:4]
  wire  success_sim_serial_out_valid; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.TinyRocketConfig.fir 209028:4]
  wire [31:0] success_sim_serial_out_bits; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.TinyRocketConfig.fir 209028:4]
  wire  success_sim_exit; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.TinyRocketConfig.fir 209028:4]
  wire  uart_sim_0_clock; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.TinyRocketConfig.fir 209044:4]
  wire  uart_sim_0_reset; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.TinyRocketConfig.fir 209044:4]
  wire  uart_sim_0_io_uart_txd; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.TinyRocketConfig.fir 209044:4]
  wire  uart_sim_0_io_uart_rxd; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.TinyRocketConfig.fir 209044:4]
  wire  dtm_success = SimJTAG_exit == 32'h1; // @[Periphery.scala 233:26 chipyard.TestHarness.TinyRocketConfig.fir 209002:4]
  wire  _T_2 = ~reset; // @[HarnessBinders.scala 190:105 chipyard.TestHarness.TinyRocketConfig.fir 208990:4]
  wire  _T_3 = SimJTAG_exit >= 32'h2; // @[Periphery.scala 234:19 chipyard.TestHarness.TinyRocketConfig.fir 209004:4]
  wire [31:0] _T_4 = {{1'd0}, SimJTAG_exit[31:1]}; // @[Periphery.scala 235:59 chipyard.TestHarness.TinyRocketConfig.fir 209006:6]
  ChipTop chiptop ( // @[TestHarness.scala 34:19 chipyard.TestHarness.TinyRocketConfig.fir 208969:4]
    .jtag_TCK(chiptop_jtag_TCK),
    .jtag_TMS(chiptop_jtag_TMS),
    .jtag_TDI(chiptop_jtag_TDI),
    .jtag_TDO_data(chiptop_jtag_TDO_data),
    .jtag_TDO_driven(chiptop_jtag_TDO_driven),
    .serial_tl_clock(chiptop_serial_tl_clock),
    .serial_tl_bits_in_ready(chiptop_serial_tl_bits_in_ready),
    .serial_tl_bits_in_valid(chiptop_serial_tl_bits_in_valid),
    .serial_tl_bits_in_bits(chiptop_serial_tl_bits_in_bits),
    .serial_tl_bits_out_ready(chiptop_serial_tl_bits_out_ready),
    .serial_tl_bits_out_valid(chiptop_serial_tl_bits_out_valid),
    .serial_tl_bits_out_bits(chiptop_serial_tl_bits_out_bits),
    .uart_0_txd(chiptop_uart_0_txd),
    .uart_0_rxd(chiptop_uart_0_rxd),
    .reset_wire_reset(chiptop_reset_wire_reset),
    .clock(chiptop_clock)
  );
  SimJTAG #(.TICK_DELAY(3)) SimJTAG ( // @[HarnessBinders.scala 190:26 chipyard.TestHarness.TinyRocketConfig.fir 208981:4]
    .clock(SimJTAG_clock),
    .reset(SimJTAG_reset),
    .jtag_TRSTn(SimJTAG_jtag_TRSTn),
    .jtag_TCK(SimJTAG_jtag_TCK),
    .jtag_TMS(SimJTAG_jtag_TMS),
    .jtag_TDI(SimJTAG_jtag_TDI),
    .jtag_TDO_data(SimJTAG_jtag_TDO_data),
    .jtag_TDO_driven(SimJTAG_jtag_TDO_driven),
    .enable(SimJTAG_enable),
    .init_done(SimJTAG_init_done),
    .exit(SimJTAG_exit)
  );
  plusarg_reader #(.FORMAT("jtag_rbb_enable=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.TinyRocketConfig.fir 208998:4]
    .out(plusarg_reader_out)
  );
  SerialRAM_inTestHarness ram ( // @[SerialAdapter.scala 27:26 chipyard.TestHarness.TinyRocketConfig.fir 209018:4]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_ser_in_ready(ram_io_ser_in_ready),
    .io_ser_in_valid(ram_io_ser_in_valid),
    .io_ser_in_bits(ram_io_ser_in_bits),
    .io_ser_out_ready(ram_io_ser_out_ready),
    .io_ser_out_valid(ram_io_ser_out_valid),
    .io_ser_out_bits(ram_io_ser_out_bits),
    .io_tsi_ser_in_ready(ram_io_tsi_ser_in_ready),
    .io_tsi_ser_in_valid(ram_io_tsi_ser_in_valid),
    .io_tsi_ser_in_bits(ram_io_tsi_ser_in_bits),
    .io_tsi_ser_out_ready(ram_io_tsi_ser_out_ready),
    .io_tsi_ser_out_valid(ram_io_tsi_ser_out_valid),
    .io_tsi_ser_out_bits(ram_io_tsi_ser_out_bits)
  );
  SimSerial success_sim ( // @[SerialAdapter.scala 37:23 chipyard.TestHarness.TinyRocketConfig.fir 209028:4]
    .clock(success_sim_clock),
    .reset(success_sim_reset),
    .serial_in_ready(success_sim_serial_in_ready),
    .serial_in_valid(success_sim_serial_in_valid),
    .serial_in_bits(success_sim_serial_in_bits),
    .serial_out_ready(success_sim_serial_out_ready),
    .serial_out_valid(success_sim_serial_out_valid),
    .serial_out_bits(success_sim_serial_out_bits),
    .exit(success_sim_exit)
  );
  UARTAdapter_inTestHarness uart_sim_0 ( // @[UARTAdapter.scala 132:28 chipyard.TestHarness.TinyRocketConfig.fir 209044:4]
    .clock(uart_sim_0_clock),
    .reset(uart_sim_0_reset),
    .io_uart_txd(uart_sim_0_io_uart_txd),
    .io_uart_rxd(uart_sim_0_io_uart_rxd)
  );
  assign io_success = success_sim_exit | dtm_success; // @[HarnessBinders.scala 236:22 chipyard.TestHarness.TinyRocketConfig.fir 209041:4 HarnessBinders.scala 236:35 chipyard.TestHarness.TinyRocketConfig.fir 209042:6]
  assign chiptop_jtag_TCK = SimJTAG_jtag_TCK; // @[Periphery.scala 220:15 chipyard.TestHarness.TinyRocketConfig.fir 208991:4]
  assign chiptop_jtag_TMS = SimJTAG_jtag_TMS; // @[Periphery.scala 221:15 chipyard.TestHarness.TinyRocketConfig.fir 208992:4]
  assign chiptop_jtag_TDI = SimJTAG_jtag_TDI; // @[Periphery.scala 222:15 chipyard.TestHarness.TinyRocketConfig.fir 208993:4]
  assign chiptop_serial_tl_bits_in_valid = ram_io_ser_in_valid; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.TinyRocketConfig.fir 209025:4]
  assign chiptop_serial_tl_bits_in_bits = ram_io_ser_in_bits; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.TinyRocketConfig.fir 209024:4]
  assign chiptop_serial_tl_bits_out_ready = ram_io_ser_out_ready; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.TinyRocketConfig.fir 209023:4]
  assign chiptop_uart_0_rxd = uart_sim_0_io_uart_rxd; // @[UARTAdapter.scala 135:18 chipyard.TestHarness.TinyRocketConfig.fir 209048:4]
  assign chiptop_reset_wire_reset = reset; // @[TestHarness.scala 41:24 chipyard.TestHarness.TinyRocketConfig.fir 208973:4]
  assign chiptop_clock = clock; // @[Clocks.scala 106:18 chipyard.TestHarness.TinyRocketConfig.fir 208975:4]
  assign SimJTAG_clock = clock; // @[Periphery.scala 225:14 chipyard.TestHarness.TinyRocketConfig.fir 208996:4]
  assign SimJTAG_reset = reset; // @[HarnessBinders.scala 190:97 chipyard.TestHarness.TinyRocketConfig.fir 208988:4]
  assign SimJTAG_jtag_TDO_data = chiptop_jtag_TDO_data; // @[Periphery.scala 223:17 chipyard.TestHarness.TinyRocketConfig.fir 208995:4]
  assign SimJTAG_jtag_TDO_driven = chiptop_jtag_TDO_driven; // @[Periphery.scala 223:17 chipyard.TestHarness.TinyRocketConfig.fir 208994:4]
  assign SimJTAG_enable = plusarg_reader_out[0]; // @[Periphery.scala 228:18 chipyard.TestHarness.TinyRocketConfig.fir 209000:4]
  assign SimJTAG_init_done = ~reset; // @[HarnessBinders.scala 190:105 chipyard.TestHarness.TinyRocketConfig.fir 208990:4]
  assign ram_clock = chiptop_serial_tl_clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 209019:4]
  assign ram_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 208971:4 chipyard.TestHarness.TinyRocketConfig.fir 208972:4]
  assign ram_io_ser_in_ready = chiptop_serial_tl_bits_in_ready; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.TinyRocketConfig.fir 209026:4]
  assign ram_io_ser_out_valid = chiptop_serial_tl_bits_out_valid; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.TinyRocketConfig.fir 209022:4]
  assign ram_io_ser_out_bits = chiptop_serial_tl_bits_out_bits; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.TinyRocketConfig.fir 209021:4]
  assign ram_io_tsi_ser_in_valid = success_sim_serial_in_valid; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.TinyRocketConfig.fir 209039:4]
  assign ram_io_tsi_ser_in_bits = success_sim_serial_in_bits; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.TinyRocketConfig.fir 209038:4]
  assign ram_io_tsi_ser_out_ready = success_sim_serial_out_ready; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.TinyRocketConfig.fir 209037:4]
  assign success_sim_clock = chiptop_serial_tl_clock; // @[SerialAdapter.scala 38:20 chipyard.TestHarness.TinyRocketConfig.fir 209033:4]
  assign success_sim_reset = reset; // @[HarnessBinders.scala 235:103 chipyard.TestHarness.TinyRocketConfig.fir 209027:4]
  assign success_sim_serial_in_ready = ram_io_tsi_ser_in_ready; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.TinyRocketConfig.fir 209040:4]
  assign success_sim_serial_out_valid = ram_io_tsi_ser_out_valid; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.TinyRocketConfig.fir 209036:4]
  assign success_sim_serial_out_bits = ram_io_tsi_ser_out_bits; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.TinyRocketConfig.fir 209035:4]
  assign uart_sim_0_clock = clock; // @[chipyard.TestHarness.TinyRocketConfig.fir 209045:4]
  assign uart_sim_0_reset = reset; // @[chipyard.TestHarness.TinyRocketConfig.fir 209046:4]
  assign uart_sim_0_io_uart_txd = chiptop_uart_0_txd; // @[UARTAdapter.scala 134:28 chipyard.TestHarness.TinyRocketConfig.fir 209047:4]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & _T_2) begin
          $fwrite(32'h80000002,"*** FAILED *** (exit code = %d)\n",_T_4); // @[Periphery.scala 235:13 chipyard.TestHarness.TinyRocketConfig.fir 209010:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3 & _T_2) begin
          $fatal; // @[Periphery.scala 236:11 chipyard.TestHarness.TinyRocketConfig.fir 209015:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module mem_inTestHarness(
  input  [9:0] RW0_addr,
  input        RW0_en,
  input        RW0_clk,
  input        RW0_wmode,
  input  [7:0] RW0_wdata_0,
  input  [7:0] RW0_wdata_1,
  input  [7:0] RW0_wdata_2,
  input  [7:0] RW0_wdata_3,
  output [7:0] RW0_rdata_0,
  output [7:0] RW0_rdata_1,
  output [7:0] RW0_rdata_2,
  output [7:0] RW0_rdata_3,
  input        RW0_wmask_0,
  input        RW0_wmask_1,
  input        RW0_wmask_2,
  input        RW0_wmask_3
);
  wire [9:0] mem_ext_RW0_addr;
  wire  mem_ext_RW0_en;
  wire  mem_ext_RW0_clk;
  wire  mem_ext_RW0_wmode;
  wire [31:0] mem_ext_RW0_wdata;
  wire [31:0] mem_ext_RW0_rdata;
  wire [3:0] mem_ext_RW0_wmask;
  wire [15:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [15:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  mem_ext mem_ext (
    .RW0_addr(mem_ext_RW0_addr),
    .RW0_en(mem_ext_RW0_en),
    .RW0_clk(mem_ext_RW0_clk),
    .RW0_wmode(mem_ext_RW0_wmode),
    .RW0_wdata(mem_ext_RW0_wdata),
    .RW0_rdata(mem_ext_RW0_rdata),
    .RW0_wmask(mem_ext_RW0_wmask)
  );
  assign mem_ext_RW0_clk = RW0_clk;
  assign mem_ext_RW0_en = RW0_en;
  assign mem_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = mem_ext_RW0_rdata[7:0];
  assign RW0_rdata_1 = mem_ext_RW0_rdata[15:8];
  assign RW0_rdata_2 = mem_ext_RW0_rdata[23:16];
  assign RW0_rdata_3 = mem_ext_RW0_rdata[31:24];
  assign mem_ext_RW0_wmode = RW0_wmode;
  assign mem_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign mem_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
